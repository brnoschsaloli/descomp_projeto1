library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Operacao_ULA_2bits, habLeituraMEM, habEscritaMEM 
      -- Inicializa os endereços:
tmp(0) := "00" & x"9" & '1' & x"B5";	-- JSR ZERA_INCREMENTO	#ZERA AS POSICOES DE MEMORIA QUE ARMAZENAM O INCREMENTO
tmp(1) := "00" & x"9" & '1' & x"AB";	-- JSR ZERA_DECREMENTO	#ZERA AS POSICOES DE MEMORIA QUE ARMAZENAM O DECREMENTO
tmp(2) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(3) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(4) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do registrador no LDR8
tmp(5) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do registrador no LDR9
tmp(6) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(7) := "00" & x"5" & '1' & x"20";	-- STA 288, R0	#ZERA HEX0
tmp(8) := "00" & x"5" & '1' & x"21";	-- STA 289, R0	#ZERA HEX1
tmp(9) := "00" & x"5" & '1' & x"22";	-- STA 290, R0	#ZERA HEX2
tmp(10) := "00" & x"5" & '1' & x"23";	-- STA 291, R0	#ZERA HEX3
tmp(11) := "00" & x"5" & '1' & x"24";	-- STA 292, R0	#ZERA HEX4
tmp(12) := "00" & x"5" & '1' & x"25";	-- STA 293, R0	#ZERA HEX5
tmp(13) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do registrador em MEM[9] (flag de decremento)
tmp(14) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega o registrador com o valor 9
tmp(15) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do registrador em MEM[10] (inibir unidade)
tmp(16) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do registrador em MEM[11] (inibir dezena)
tmp(17) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do registrador em MEM[12] (inibir centena)
tmp(18) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do registrador em MEM[13] (inibir milhar)
tmp(19) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do registrador em MEM[14] (inibir dezena de milhar)
tmp(20) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do registrador em MEM[15] (inibir centena de milhar)
tmp(21) := "11" & x"4" & '0' & x"08";	-- LDI 8, R3	#COLUNA 8
tmp(22) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(23) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(24) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(25) := "11" & x"4" & '0' & x"3A";	-- LDI 58, R3	#dois pontos
tmp(26) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(27) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(28) := "11" & x"4" & '0' & x"0B";	-- LDI 11, R3	#COLUNA 11
tmp(29) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(30) := "11" & x"4" & '0' & x"3A";	-- LDI 58, R3	#dois pontos
tmp(31) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(32) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(33) := "00" & x"1" & '0' & x"09";	-- LDA 9, R0	#Carrega o registrador com a leitura de MEM[9] (flag de decremento)
tmp(34) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(35) := "00" & x"7" & '0' & x"2B";	-- JEQ FLAG_DESATIVADA	#Desvia se igual a 0 (botão não foi pressionado)
tmp(36) := "00" & x"1" & '1' & x"62";	-- LDA 354, R0	#Carrega o registrador com a leitura do botão KEY2
tmp(37) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(38) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(39) := "00" & x"7" & '0' & x"30";	-- JEQ NAO_CLICOU0	#Desvia se igual a 0 (botão não foi pressionado)
tmp(40) := "00" & x"9" & '1' & x"68";	-- JSR DECREMENTO
tmp(41) := "00" & x"9" & '0' & x"42";	-- JSR INCREMENTO	#O botão foi pressionado, chama a sub-rotina de decremento
tmp(42) := "00" & x"6" & '0' & x"30";	-- JMP NAO_CLICOU0
tmp(43) := "00" & x"1" & '1' & x"60";	-- LDA 352, R0	#Carrega o registrador com a leitura do botão KEY0
tmp(44) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(45) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(46) := "00" & x"7" & '0' & x"30";	-- JEQ NAO_CLICOU0	#Desvia se igual a 0 (botão não foi pressionado)
tmp(47) := "00" & x"9" & '0' & x"42";	-- JSR INCREMENTO	#O botão foi pressionado, chama a sub-rotina de incremento
tmp(48) := "00" & x"9" & '0' & x"8D";	-- JSR SALVA_DISP	#Escreve o valor das váriaveis de contagem nos displays
tmp(49) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o registrador com a leitura do botão KEY1
tmp(50) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(51) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(52) := "00" & x"7" & '0' & x"36";	-- JEQ NAO_CLICOU1	#Desvia se igual a 0 (botão não foi pressionado)
tmp(53) := "00" & x"9" & '1' & x"28";	-- JSR DEFINE_LIM	#O botão foi pressionado, chama a sub-rotina de definir limite
tmp(54) := "00" & x"9" & '1' & x"04";	-- JSR VERIFICA_LIM
tmp(55) := "00" & x"1" & '1' & x"63";	-- LDA 355, R0	#Carrega o registrador com a leitura do botão KEY3
tmp(56) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(57) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(58) := "00" & x"7" & '0' & x"3C";	-- JEQ NAO_CLICOU2	#Desvia se igual a 0 (botão não foi pressionado)
tmp(59) := "00" & x"9" & '1' & x"C8";	-- JSR TEMPORIZADOR	#O botão foi pressionado, chama a sub-rotina de temporizador
tmp(60) := "00" & x"1" & '1' & x"64";	-- LDA 356, R0	#Carrega o registrador com a leitura do botão FPGA_RESET
tmp(61) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(62) := "00" & x"D" & '0' & x"01";	-- CEQi 1, R0	#Compara com constante 1
tmp(63) := "00" & x"7" & '0' & x"41";	-- JEQ REINICIO	#Desvia se igual a 1 (botão não foi pressionado)
tmp(64) := "00" & x"9" & '0' & x"EA";	-- JSR RESET	#O botão foi pressionado, chama a sub-rotina de reset
tmp(65) := "00" & x"6" & '0' & x"21";	-- JMP INICIO	#Fecha o laço principal, faz uma nova leitura de KEY0
tmp(66) := "10" & x"1" & '1' & x"42";	-- LDA 322, R2	#Carrega valor de SW9 no registrador 2
tmp(67) := "10" & x"5" & '1' & x"02";	-- STA 258, R2	#Escreve o valor de R2 no LED9
tmp(68) := "00" & x"5" & '1' & x"FF";	-- STA 511, R0	#Limpa a leitura do botão
tmp(69) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	#Carrega o valor de MEM[0] (contador)
tmp(70) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(71) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(72) := "00" & x"7" & '0' & x"4B";	-- JEQ VAIUM_D	#Realiza o carry out caso valor igual a 10
tmp(73) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Salva o incremento em MEM[0] (contador)
tmp(74) := "00" & x"A" & '0' & x"00";	-- RET	#Retorna da sub-rotina
tmp(75) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no registrador 0
tmp(76) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do registrador em MEM[0] (unidades)
tmp(77) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	#Carrega valor de MEM[1] no registrador (dezenas)
tmp(78) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(79) := "00" & x"D" & '0' & x"06";	-- CEQi 6, R0	#Compara o valor com constante 10
tmp(80) := "00" & x"7" & '0' & x"53";	-- JEQ VAIUM_C	#Realiza o carry out caso valor igual a 10
tmp(81) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Salva o incremento em MEM[1] (dezenas)
tmp(82) := "00" & x"A" & '0' & x"00";	-- RET
tmp(83) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no registrador
tmp(84) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do registrador em MEM[1] (dezenas)
tmp(85) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	#Carrega valor de MEM[2] no registrador (centenas)
tmp(86) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(87) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(88) := "00" & x"7" & '0' & x"5B";	-- JEQ VAIUM_M	#Realiza o carry out caso valor igual a 10
tmp(89) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Salva o incremento em MEM[2] (centenas)
tmp(90) := "00" & x"A" & '0' & x"00";	-- RET
tmp(91) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no registrador
tmp(92) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do registrador em MEM[2] (centenas)
tmp(93) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	#Carrega valor de MEM[6] no registrador (milhares)
tmp(94) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(95) := "00" & x"D" & '0' & x"06";	-- CEQi 6, R0	#Compara o valor com constante 10
tmp(96) := "00" & x"7" & '0' & x"63";	-- JEQ VAIUM_DM	#Realiza o carry out caso valor igual a 10
tmp(97) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Salva o incremento em MEM[6] (milhares)
tmp(98) := "00" & x"A" & '0' & x"00";	-- RET
tmp(99) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no registrador
tmp(100) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do registrador em MEM[6] (milhares)
tmp(101) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	#Carrega valor de MEM[7] no registrador (dezenas de milhares)
tmp(102) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(103) := "01" & x"1" & '0' & x"08";	-- LDA 8, R1	#Carrega valor de MEM[8] no registrador (centenas de milhares)
tmp(104) := "10" & x"1" & '1' & x"42";	-- LDA 322, R2	#Carrega valor de SW9 no registrador 2
tmp(105) := "10" & x"D" & '0' & x"00";	-- CEQi 0, R2	#Compara o valor do R2 com constante 0 (verifica se a chave am pm esta ligada)
tmp(106) := "00" & x"7" & '0' & x"7C";	-- JEQ 24HORAS
tmp(107) := "01" & x"D" & '0' & x"01";	-- CEQi 1, R1	#Compara o valor com constante 1
tmp(108) := "00" & x"7" & '0' & x"70";	-- JEQ COMPARA3	#Pula para o fim da rotina
tmp(109) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(110) := "00" & x"7" & '0' & x"74";	-- JEQ VAIUM_CM2	#Realiza o carry out caso valor igual a 10
tmp(111) := "00" & x"6" & '0' & x"83";	-- JMP END_DM
tmp(112) := "00" & x"D" & '0' & x"03";	-- CEQi 3, R0	#Compara o valor com constante 3
tmp(113) := "00" & x"7" & '0' & x"74";	-- JEQ VAIUM_CM2	#Realiza o carry out caso valor igual a 3
tmp(114) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Salva o incremento em MEM[7] (dezenas de milhares)
tmp(115) := "00" & x"A" & '0' & x"00";	-- RET
tmp(116) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no registrador
tmp(117) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do registrador em MEM[7] (dezenas milhares)
tmp(118) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega valor de MEM[8] no registrador (centenas de milhares)
tmp(119) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(120) := "00" & x"D" & '0' & x"02";	-- CEQi 2, R0	#Compara o valor com constante 3
tmp(121) := "00" & x"7" & '1' & x"BF";	-- JEQ ZERA_HEX_AM	#Zera se chegar ao final
tmp(122) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Salva o incremento em MEM[8] (centena de milhares)
tmp(123) := "00" & x"A" & '0' & x"00";	-- RET
tmp(124) := "01" & x"D" & '0' & x"02";	-- CEQi 2, R1	#Compara o valor com constante 2
tmp(125) := "00" & x"7" & '0' & x"81";	-- JEQ COMPARA4	#Pula para o fim da rotina
tmp(126) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(127) := "00" & x"7" & '0' & x"85";	-- JEQ VAIUM_CM	#Realiza o carry out caso valor igual a 10
tmp(128) := "00" & x"6" & '0' & x"83";	-- JMP END_DM
tmp(129) := "00" & x"D" & '0' & x"04";	-- CEQi 4, R0	#Compara o valor com constante 4
tmp(130) := "00" & x"7" & '0' & x"85";	-- JEQ VAIUM_CM	#Realiza o carry out caso valor igual a 4
tmp(131) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Salva o incremento em MEM[7] (dezenas de milhares)
tmp(132) := "00" & x"A" & '0' & x"00";	-- RET
tmp(133) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no registrador
tmp(134) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do registrador em MEM[7] (dezenas milhares)
tmp(135) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega valor de MEM[8] no registrador (centenas de milhares)
tmp(136) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(137) := "00" & x"D" & '0' & x"03";	-- CEQi 3, R0	#Compara o valor com constante 3
tmp(138) := "00" & x"7" & '1' & x"B5";	-- JEQ ZERA_INCREMENTO	#Zera se chegar ao final
tmp(139) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Salva o incremento em MEM[8] (centena de milhares)
tmp(140) := "00" & x"A" & '0' & x"00";	-- RET
tmp(141) := "00" & x"1" & '0' & x"09";	-- LDA 9, R0
tmp(142) := "00" & x"D" & '0' & x"01";	-- CEQi 1, R0
tmp(143) := "00" & x"7" & '0' & x"BD";	-- JEQ SALVA_DECREMENTO
tmp(144) := "11" & x"4" & '0' & x"0D";	-- LDI 13, R3	#COLUNA 13
tmp(145) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(146) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(147) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(148) := "11" & x"1" & '0' & x"00";	-- LDA 0, R3	#Carrega o valor de MEM[0] (unidades)
tmp(149) := "11" & x"5" & '1' & x"20";	-- STA 288, R3	#Armazena valor do registrador de unidades no HEX0
tmp(150) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(151) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(152) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(153) := "11" & x"4" & '0' & x"0C";	-- LDI 12, R3	#COLUNA 12
tmp(154) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(155) := "11" & x"1" & '0' & x"01";	-- LDA 1, R3	#Carrega o valor de MEM[1] (dezenas)
tmp(156) := "11" & x"5" & '1' & x"21";	-- STA 289, R3	#Armazena valor do registrador de dezenas no HEX1
tmp(157) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(158) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(159) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(160) := "11" & x"4" & '0' & x"0A";	-- LDI 10, R3	#COLUNA 10
tmp(161) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(162) := "11" & x"1" & '0' & x"02";	-- LDA 2, R3	#Carrega o valor de MEM[2] (centenas)
tmp(163) := "11" & x"5" & '1' & x"22";	-- STA 290, R3	#Armazena valor do registrador de centenas no HEX2
tmp(164) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(165) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(166) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(167) := "11" & x"4" & '0' & x"09";	-- LDI 9, R3	#COLUNA 9
tmp(168) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(169) := "11" & x"1" & '0' & x"06";	-- LDA 6, R3	#Carrega o valor de MEM[6] (milhares)
tmp(170) := "11" & x"5" & '1' & x"23";	-- STA 291, R3	#Armazena valor do registrador de unidades no HEX3
tmp(171) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(172) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(173) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(174) := "11" & x"4" & '0' & x"07";	-- LDI 7, R3	#COLUNA 7
tmp(175) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(176) := "11" & x"1" & '0' & x"07";	-- LDA 7, R3	#Carrega o valor de MEM[7] (dezenas de milhares)
tmp(177) := "11" & x"5" & '1' & x"24";	-- STA 292, R3	#Armazena valor do registrador de dezenas no HEX4
tmp(178) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(179) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(180) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(181) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#COLUNA 6
tmp(182) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(183) := "11" & x"1" & '0' & x"08";	-- LDA 8, R3	#Carrega o valor de MEM[8] (centenas de milhares)
tmp(184) := "11" & x"5" & '1' & x"25";	-- STA 293, R3	#Armazena valor do registrador de centenas no HEX5
tmp(185) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(186) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(187) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(188) := "00" & x"A" & '0' & x"00";	-- RET
tmp(189) := "11" & x"4" & '0' & x"0D";	-- LDI 13, R3	#COLUNA 13
tmp(190) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(191) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(192) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(193) := "11" & x"1" & '0' & x"1E";	-- LDA 30, R3	#Carrega o valor de MEM[30] (unidades)
tmp(194) := "11" & x"5" & '1' & x"20";	-- STA 288, R3	#Armazena valor do registrador de unidades no HEX0
tmp(195) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(196) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(197) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(198) := "11" & x"4" & '0' & x"0C";	-- LDI 12, R3	#COLUNA 12
tmp(199) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(200) := "11" & x"1" & '0' & x"1F";	-- LDA 31, R3	#Carrega o valor de MEM[31] (dezenas)
tmp(201) := "11" & x"5" & '1' & x"21";	-- STA 289, R3	#Armazena valor do registrador de dezenas no HEX1
tmp(202) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(203) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(204) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(205) := "11" & x"4" & '0' & x"0A";	-- LDI 10, R3	#COLUNA 10
tmp(206) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(207) := "11" & x"1" & '0' & x"20";	-- LDA 32, R3	#Carrega o valor de MEM[32] (centenas)
tmp(208) := "11" & x"5" & '1' & x"22";	-- STA 290, R3	#Armazena valor do registrador de centenas no HEX2
tmp(209) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(210) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(211) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(212) := "11" & x"4" & '0' & x"09";	-- LDI 9, R3	#COLUNA 9
tmp(213) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(214) := "11" & x"1" & '0' & x"21";	-- LDA 33, R3	#Carrega o valor de MEM[33] (milhares)
tmp(215) := "11" & x"5" & '1' & x"23";	-- STA 291, R3	#Armazena valor do registrador de unidades no HEX3
tmp(216) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(217) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(218) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(219) := "11" & x"4" & '0' & x"07";	-- LDI 7, R3	#COLUNA 7
tmp(220) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(221) := "11" & x"1" & '0' & x"22";	-- LDA 34, R3	#Carrega o valor de MEM[34] (dezenas de milhares)
tmp(222) := "11" & x"5" & '1' & x"24";	-- STA 292, R3	#Armazena valor do registrador de dezenas no HEX4
tmp(223) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(224) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(225) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(226) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#COLUNA 6
tmp(227) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(228) := "11" & x"1" & '0' & x"23";	-- LDA 35, R3	#Carrega o valor de MEM[35] (centenas de milhares)
tmp(229) := "11" & x"5" & '1' & x"25";	-- STA 293, R3	#Armazena valor do registrador de centenas no HEX5
tmp(230) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(231) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(232) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(233) := "00" & x"A" & '0' & x"00";	-- RET
tmp(234) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(235) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do registrador na MEM[0] (unidades)
tmp(236) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do registrador na MEM[1] (dezenas)
tmp(237) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do registrador na MEM[2] (centenas)
tmp(238) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do registrador na MEM[6] (milhar)
tmp(239) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do registrador na MEM[7] (dezena de milhar)
tmp(240) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do registrador na MEM[8] (centena de milhar)
tmp(241) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do registrador na MEM[9] (flag de decremento)
tmp(242) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do registrador no LDR8
tmp(243) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega o registrador com o valor 9
tmp(244) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do registrador em MEM[10] (inibir unidade)
tmp(245) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do registrador em MEM[11] (inibir dezena)
tmp(246) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do registrador em MEM[12] (inibir centena)
tmp(247) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do registrador em MEM[13] (inibir milhar)
tmp(248) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do registrador em MEM[14] (inibir dezena de milhar)
tmp(249) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do registrador em MEM[15] (inibir centena de milhar)
tmp(250) := "11" & x"4" & '0' & x"0A";	-- LDI 10, R3	#COLUNA 10
tmp(251) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(252) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#LINHA 6
tmp(253) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(254) := "11" & x"4" & '0' & x"00";	-- LDI 0, R3	#zera o sino
tmp(255) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(256) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(257) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(258) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(259) := "00" & x"A" & '0' & x"00";	-- RET
tmp(260) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	#Carrega o valor de MEM[0] (unidades)
tmp(261) := "00" & x"8" & '0' & x"0A";	-- CEQ 10, R0	#Compara o valor de MEM[10] (inibir unidade)
tmp(262) := "00" & x"7" & '1' & x"08";	-- JEQ NEXT_LIM1
tmp(263) := "00" & x"A" & '0' & x"00";	-- RET
tmp(264) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	#Carrega o valor de MEM[1] (dezenas)
tmp(265) := "00" & x"8" & '0' & x"0B";	-- CEQ 11, R0	#Compara o valor de MEM[11] (inibir dezenas)
tmp(266) := "00" & x"7" & '1' & x"0C";	-- JEQ NEXT_LIM2
tmp(267) := "00" & x"A" & '0' & x"00";	-- RET
tmp(268) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	#Carrega o valor de MEM[2] (centenas)
tmp(269) := "00" & x"8" & '0' & x"0C";	-- CEQ 12, R0	#Compara o valor de MEM[12] (inibir centenas)
tmp(270) := "00" & x"7" & '1' & x"10";	-- JEQ NEXT_LIM3
tmp(271) := "00" & x"A" & '0' & x"00";	-- RET
tmp(272) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	#Carrega o valor de MEM[6] (milhar)
tmp(273) := "00" & x"8" & '0' & x"0D";	-- CEQ 13, R0	#Compara o valor de MEM[13] (inibir milhar)
tmp(274) := "00" & x"7" & '1' & x"14";	-- JEQ NEXT_LIM4
tmp(275) := "00" & x"A" & '0' & x"00";	-- RET
tmp(276) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	#Carrega o valor de MEM[7] (dezena de milhar)
tmp(277) := "00" & x"8" & '0' & x"0E";	-- CEQ 14, R0	#Compara o valor de MEM[10] (inibir dezena de milhar)
tmp(278) := "00" & x"7" & '1' & x"18";	-- JEQ NEXT_LIM5
tmp(279) := "00" & x"A" & '0' & x"00";	-- RET
tmp(280) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega o valor de MEM[8] (centena de milhar)
tmp(281) := "00" & x"8" & '0' & x"0F";	-- CEQ 15, R0	#Compara o valor de MEM[10] (inibir centena de milhar)
tmp(282) := "00" & x"7" & '1' & x"1C";	-- JEQ TODOS_IGUAL
tmp(283) := "00" & x"A" & '0' & x"00";	-- RET
tmp(284) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o registrador com o valor 1
tmp(285) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do registrador no LDR8
tmp(286) := "11" & x"4" & '0' & x"0A";	-- LDI 10, R3	#COLUNA 10
tmp(287) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(288) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#LINHA 6
tmp(289) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(290) := "11" & x"4" & '0' & x"1F";	-- LDI 31, R3	#sino
tmp(291) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(292) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(293) := "00" & x"4" & '0' & x"FF";	-- LDI 255, R0	#Carrega o registrador com o valor 255
tmp(294) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(295) := "00" & x"A" & '0' & x"00";	-- RET
tmp(296) := "11" & x"4" & '0' & x"0A";	-- LDI 10, R3	#COLUNA 10
tmp(297) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(298) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#LINHA 6
tmp(299) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(300) := "11" & x"4" & '0' & x"00";	-- LDI 0, R3	#zera o sino
tmp(301) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(302) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(303) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(304) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(305) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(306) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do registrador no LDR8
tmp(307) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(308) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(309) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do registrador em MEM[10] (inibir unidade)
tmp(310) := "00" & x"4" & '0' & x"04";	-- LDI 4, R0	#Carrega o registrador com o valor 4
tmp(311) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(312) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o registrador com a leitura do botão KEY1
tmp(313) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(314) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(315) := "00" & x"7" & '1' & x"38";	-- JEQ AGUARDA_D	#Desvia se igual a 0 (botão não foi pressionado)
tmp(316) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(317) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(318) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do registrador em MEM[11] (inibir dezena)
tmp(319) := "00" & x"4" & '0' & x"10";	-- LDI 16, R0	#Carrega o registrador com o valor 16
tmp(320) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(321) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o registrador com a leitura do botão KEY1
tmp(322) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(323) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(324) := "00" & x"7" & '1' & x"41";	-- JEQ AGUARDA_C	#Desvia se igual a 0 (botão não foi pressionado)
tmp(325) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(326) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(327) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do registrador em MEM[12] (inibir centena)
tmp(328) := "00" & x"4" & '0' & x"20";	-- LDI 32, R0	#Carrega o registrador com o valor 32
tmp(329) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(330) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o registrador com a leitura do botão KEY1
tmp(331) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(332) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(333) := "00" & x"7" & '1' & x"4A";	-- JEQ AGUARDA_M	#Desvia se igual a 0 (botão não foi pressionado)
tmp(334) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(335) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(336) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do registrador em MEM[13] (inibir milhar)
tmp(337) := "00" & x"4" & '0' & x"80";	-- LDI 128, R0	#Carrega o registrador com o valor 128
tmp(338) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(339) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o registrador com a leitura do botão KEY1
tmp(340) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(341) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(342) := "00" & x"7" & '1' & x"53";	-- JEQ AGUARDA_DM	#Desvia se igual a 0 (botão não foi pressionado)
tmp(343) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(344) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(345) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do registrador em MEM[13] (inibir dezena de milhar)
tmp(346) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(347) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(348) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o registrador com o valor 1
tmp(349) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do registrador no LDR9
tmp(350) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o registrador com a leitura do botão KEY1
tmp(351) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(352) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(353) := "00" & x"7" & '1' & x"5E";	-- JEQ AGUARDA_CM	#Desvia se igual a 0 (botão não foi pressionado)
tmp(354) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(355) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(356) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do registrador em MEM[15] (inibir centena de milhar)
tmp(357) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(358) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do registrador no LDR9
tmp(359) := "00" & x"A" & '0' & x"00";	-- RET
tmp(360) := "11" & x"4" & '0' & x"0A";	-- LDI 10, R3	#COLUNA 10
tmp(361) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(362) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#LINHA 6
tmp(363) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(364) := "11" & x"4" & '0' & x"00";	-- LDI 0, R3	#zera o sino
tmp(365) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(366) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(367) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(368) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(369) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega 0 para o registrador
tmp(370) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do registrador no LDR8
tmp(371) := "00" & x"5" & '1' & x"FD";	-- STA 509, R0	#Limpa a leitura do botão KEY2
tmp(372) := "00" & x"1" & '0' & x"1E";	-- LDA 30, R0	#Carrega MEM[30] (unidades decremento) no registrador
tmp(373) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Verifica se MEM[30] == 0
tmp(374) := "00" & x"7" & '1' & x"7A";	-- JEQ VEMUM_D	#Se MEM[30] == 0, realiza o "empréstimo"
tmp(375) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	#Subtrai 1 de MEM[0]
tmp(376) := "00" & x"5" & '0' & x"1E";	-- STA 30, R0	#Armazena o novo valor de MEM[30]
tmp(377) := "00" & x"A" & '0' & x"00";	-- RET	#Retorna da sub-rotina
tmp(378) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega 9 no registrador
tmp(379) := "00" & x"5" & '0' & x"1E";	-- STA 30, R0	#Define MEM[30] para 9
tmp(380) := "00" & x"1" & '0' & x"1F";	-- LDA 31, R0	#Carrega MEM[31] (dezenas decremento) no registrador
tmp(381) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Verifica se MEM[1] == 0
tmp(382) := "00" & x"7" & '1' & x"82";	-- JEQ VEMUM_C	#Se MEM[31] == 0, realiza o próximo "empréstimo"
tmp(383) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	#Subtrai 1 de MEM[1]
tmp(384) := "00" & x"5" & '0' & x"1F";	-- STA 31, R0	#Armazena o novo valor de MEM[31]
tmp(385) := "00" & x"A" & '0' & x"00";	-- RET	#Retorna da sub-rotina
tmp(386) := "00" & x"4" & '0' & x"05";	-- LDI 5, R0	#Carrega 5 no registrador
tmp(387) := "00" & x"5" & '0' & x"1F";	-- STA 31, R0	#Define MEM[31] para 5
tmp(388) := "00" & x"1" & '0' & x"20";	-- LDA 32, R0	#Carrega MEM[32] (centenas decremento) no registrador
tmp(389) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Verifica se MEM[2] == 0
tmp(390) := "00" & x"7" & '1' & x"8A";	-- JEQ VEMUM_M	#Se MEM[32] == 0, realiza o próximo "empréstimo"
tmp(391) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	#Subtrai 1 de MEM[2]
tmp(392) := "00" & x"5" & '0' & x"20";	-- STA 32, R0	#Armazena o novo valor de MEM[32]
tmp(393) := "00" & x"A" & '0' & x"00";	-- RET	#Retorna da sub-rotina
tmp(394) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega 9 no registrador
tmp(395) := "00" & x"5" & '0' & x"20";	-- STA 32, R0	#Define MEM[32] para 9
tmp(396) := "00" & x"1" & '0' & x"21";	-- LDA 33, R0	#Carrega MEM[33] (milhares decremento) no registrador
tmp(397) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Verifica se MEM[33] == 0
tmp(398) := "00" & x"7" & '1' & x"92";	-- JEQ VEMUM_DM	#Se MEM[33] == 0, realiza o próximo "empréstimo"
tmp(399) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	#Subtrai 1 de MEM[33]
tmp(400) := "00" & x"5" & '0' & x"21";	-- STA 33, R0	#Armazena o novo valor de MEM[33]
tmp(401) := "00" & x"A" & '0' & x"00";	-- RET	#Retorna da sub-rotina
tmp(402) := "00" & x"4" & '0' & x"05";	-- LDI 5, R0	#Carrega 5 no registrador
tmp(403) := "00" & x"5" & '0' & x"21";	-- STA 33, R0	#Define MEM[33] para 5
tmp(404) := "00" & x"1" & '0' & x"22";	-- LDA 34, R0	#Carrega MEM[34] (dezenas de milhares decremento) no registrador
tmp(405) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Verifica se MEM[34] == 0
tmp(406) := "00" & x"7" & '1' & x"9A";	-- JEQ VEMUM_CM	#Se MEM[34] == 0, realiza o próximo "empréstimo"
tmp(407) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	#Subtrai 1 de MEM[34]
tmp(408) := "00" & x"5" & '0' & x"22";	-- STA 34, R0	#Armazena o novo valor de MEM[34]
tmp(409) := "00" & x"A" & '0' & x"00";	-- RET	#Retorna da sub-rotina
tmp(410) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega 9 no registrador
tmp(411) := "00" & x"5" & '0' & x"22";	-- STA 34, R0	#Define MEM[34] para 9
tmp(412) := "00" & x"1" & '0' & x"23";	-- LDA 35, R0	#Carrega MEM[35] (centenas de milhares decremento) no registrador
tmp(413) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Verifica se MEM[35] == 0
tmp(414) := "11" & x"4" & '0' & x"0A";	-- LDI 10, R3	#COLUNA 10
tmp(415) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(416) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#LINHA 6
tmp(417) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(418) := "11" & x"4" & '0' & x"1F";	-- LDI 31, R3	#sino
tmp(419) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(420) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(421) := "00" & x"4" & '0' & x"FF";	-- LDI 255, R0	#Carrega o registrador com o valor 255
tmp(422) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(423) := "00" & x"7" & '1' & x"AB";	-- JEQ ZERA_DECREMENTO	#Zera se for igual a 0
tmp(424) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	#Subtrai 1 de MEM[35]
tmp(425) := "00" & x"5" & '0' & x"23";	-- STA 35, R0	#Armazena o novo valor de MEM[35]
tmp(426) := "00" & x"A" & '0' & x"00";	-- RET	#Retorna da sub-rotina
tmp(427) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(428) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do registrador no LDR9
tmp(429) := "00" & x"5" & '0' & x"1E";	-- STA 30, R0	#Armazena o valor do registrador na MEM[30] (unidades)
tmp(430) := "00" & x"5" & '0' & x"1F";	-- STA 31, R0	#Armazena o valor do registrador na MEM[31] (dezenas)
tmp(431) := "00" & x"5" & '0' & x"20";	-- STA 32, R0	#Armazena o valor do registrador na MEM[32] (centenas)
tmp(432) := "00" & x"5" & '0' & x"21";	-- STA 33, R0	#Armazena o valor do registrador na MEM[33] (milhar)
tmp(433) := "00" & x"5" & '0' & x"22";	-- STA 34, R0	#Armazena o valor do registrador na MEM[34] (dezena de milhar)
tmp(434) := "00" & x"5" & '0' & x"23";	-- STA 35, R0	#Armazena o valor do registrador na MEM[35] (centena de milhar)
tmp(435) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do registrador na MEM[9] (flag de decremento)
tmp(436) := "00" & x"A" & '0' & x"00";	-- RET
tmp(437) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(438) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do registrador no LDR9
tmp(439) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do registrador na MEM[0] (unidades)
tmp(440) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do registrador na MEM[1] (dezenas)
tmp(441) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do registrador na MEM[2] (centenas)
tmp(442) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do registrador na MEM[6] (milhar)
tmp(443) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do registrador na MEM[7] (dezena de milhar)
tmp(444) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do registrador na MEM[8] (centena de milhar)
tmp(445) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do registrador na MEM[9] (flag de decremento)
tmp(446) := "00" & x"A" & '0' & x"00";	-- RET
tmp(447) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(448) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do registrador na MEM[0] (unidades)
tmp(449) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do registrador na MEM[1] (dezenas)
tmp(450) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do registrador na MEM[2] (centenas)
tmp(451) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do registrador na MEM[6] (milhar)
tmp(452) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do registrador na MEM[8] (centena de milhar)
tmp(453) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o registrador com o valor 1
tmp(454) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do registrador na MEM[7] (dezena de milhar)
tmp(455) := "00" & x"A" & '0' & x"00";	-- RET
tmp(456) := "00" & x"5" & '1' & x"FC";	-- STA 508, R0	#Limpa a leitura do botão tres
tmp(457) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(458) := "00" & x"5" & '0' & x"1E";	-- STA 30, R0	#Armazena o valor do registrador em MEM[30] (unidade decremento)
tmp(459) := "00" & x"4" & '0' & x"04";	-- LDI 4, R0	#Carrega o registrador com o valor 4
tmp(460) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(461) := "00" & x"1" & '1' & x"63";	-- LDA 355, R0	#Carrega o registrador com a leitura do botão KEY3
tmp(462) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(463) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(464) := "00" & x"7" & '1' & x"CD";	-- JEQ AGUARDA_DT	#Desvia se igual a 0 (botão não foi pressionado)
tmp(465) := "00" & x"5" & '1' & x"FC";	-- STA 508, R0	#Limpa a leitura do botão tres
tmp(466) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(467) := "00" & x"5" & '0' & x"1F";	-- STA 31, R0	#Armazena o valor do registrador em MEM[31] (dezena decremento)
tmp(468) := "00" & x"4" & '0' & x"10";	-- LDI 16, R0	#Carrega o registrador com o valor 16
tmp(469) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(470) := "00" & x"1" & '1' & x"63";	-- LDA 355, R0	#Carrega o registrador com a leitura do botão KEY3
tmp(471) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(472) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(473) := "00" & x"7" & '1' & x"D6";	-- JEQ AGUARDA_CT	#Desvia se igual a 0 (botão não foi pressionado)
tmp(474) := "00" & x"5" & '1' & x"FC";	-- STA 508, R0	#Limpa a leitura do botão tres
tmp(475) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(476) := "00" & x"5" & '0' & x"20";	-- STA 32, R0	#Armazena o valor do registrador em MEM[32] (centena decremento)
tmp(477) := "00" & x"4" & '0' & x"20";	-- LDI 32, R0	#Carrega o registrador com o valor 32
tmp(478) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(479) := "00" & x"1" & '1' & x"63";	-- LDA 355, R0	#Carrega o registrador com a leitura do botão KEY3
tmp(480) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(481) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(482) := "00" & x"7" & '1' & x"DF";	-- JEQ AGUARDA_MT	#Desvia se igual a 0 (botão não foi pressionado)
tmp(483) := "00" & x"5" & '1' & x"FC";	-- STA 508, R0	#Limpa a leitura do botão tres
tmp(484) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(485) := "00" & x"5" & '0' & x"21";	-- STA 33, R0	#Armazena o valor do registrador em MEM[33] (unidade de milhar decremento)
tmp(486) := "00" & x"4" & '0' & x"80";	-- LDI 128, R0	#Carrega o registrador com o valor 128
tmp(487) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(488) := "00" & x"1" & '1' & x"63";	-- LDA 355, R0	#Carrega o registrador com a leitura do botão KEY3
tmp(489) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(490) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(491) := "00" & x"7" & '1' & x"E8";	-- JEQ AGUARDA_DMT	#Desvia se igual a 0 (botão não foi pressionado)
tmp(492) := "00" & x"5" & '1' & x"FC";	-- STA 508, R0	#Limpa a leitura do botão tres
tmp(493) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(494) := "00" & x"5" & '0' & x"22";	-- STA 34, R0	#Armazena o valor do registrador em MEM[34] (dezena de milhar decremento)
tmp(495) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(496) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do registrador no LDR0 ~ LEDR7
tmp(497) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o registrador com o valor 1
tmp(498) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do registrador no LDR9
tmp(499) := "00" & x"1" & '1' & x"63";	-- LDA 355, R0	#Carrega o registrador com a leitura do botão KEY3
tmp(500) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(501) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(502) := "00" & x"7" & '1' & x"F3";	-- JEQ AGUARDA_CMT	#Desvia se igual a 0 (botão não foi pressionado)
tmp(503) := "00" & x"5" & '1' & x"FC";	-- STA 508, R0	#Limpa a leitura do botão tres
tmp(504) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o registrador com a leitura do SW7TO0
tmp(505) := "00" & x"5" & '0' & x"23";	-- STA 35, R0	#Armazena o valor do registrador em MEM[35] (centena de milhar decremento)
tmp(506) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o registrador com o valor 0
tmp(507) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do registrador no LDR9
tmp(508) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o registrador com o valor 1
tmp(509) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do registrador no MEM[9] (flag de decremento)
tmp(510) := "00" & x"A" & '0' & x"00";	-- RET
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;