library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Operacao_ULA_2bits, habLeituraMEM, habEscritaMEM 
      -- Inicializa os endereços:
tmp(0) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(1) := "00" & x"5" & '1' & x"20";	-- STA 288, R0	#Armazena o valor do acumulador em HEX0
tmp(2) := "00" & x"5" & '1' & x"21";	-- STA 289, R0	#Armazena o valor do acumulador em HEX1
tmp(3) := "00" & x"5" & '1' & x"22";	-- STA 290, R0	#Armazena o valor do acumulador em HEX2
tmp(4) := "00" & x"5" & '1' & x"23";	-- STA 291, R0	#Armazena o valor do acumulador em HEX3
tmp(5) := "00" & x"5" & '1' & x"24";	-- STA 292, R0	#Armazena o valor do acumulador em HEX4
tmp(6) := "00" & x"5" & '1' & x"25";	-- STA 293, R0	#Armazena o valor do acumulador em HEX5
tmp(7) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(8) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(9) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(10) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(11) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do acumulador no LDR9
tmp(12) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(13) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(14) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador em MEM[0] (unidades)
tmp(15) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador em MEM[1] (dezenas)
tmp(16) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador em MEM[2] (centenas)
tmp(17) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador em MEM[6] (milhares)
tmp(18) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador em MEM[7] (dezenas de milhares)
tmp(19) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do acumulador em MEM[8] (centenas de milhares)
tmp(20) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador em MEM[9] (flag inibir contagem)
tmp(21) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega o acumulador com o valor 9
tmp(22) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do acumulador em MEM[10] (inibir unidade)
tmp(23) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do acumulador em MEM[11] (inibir dezena)
tmp(24) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do acumulador em MEM[12] (inibir centena)
tmp(25) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do acumulador em MEM[13] (inibir milhar)
tmp(26) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do acumulador em MEM[14] (inibir dezena de milhar)
tmp(27) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do acumulador em MEM[15] (inibir centena de milhar)
tmp(28) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(29) := "00" & x"5" & '1' & x"FF";	-- STA 511, R0	#Limpa a leitura do botão zero
tmp(30) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(31) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(32) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(33) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(34) := "11" & x"4" & '0' & x"03";	-- LDI 3, R3	#COLUNA 3
tmp(35) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(36) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(37) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(38) := "11" & x"4" & '0' & x"12";	-- LDI 18, R3	#R
tmp(39) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(40) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(41) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#COLUNA 4
tmp(42) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(43) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(44) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(45) := "11" & x"4" & '0' & x"05";	-- LDI 5, R3	#E
tmp(46) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(47) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(48) := "11" & x"4" & '0' & x"05";	-- LDI 5, R3	#COLUNA 5
tmp(49) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(50) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(51) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(52) := "11" & x"4" & '0' & x"0C";	-- LDI 12, R3	#L
tmp(53) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(54) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(55) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#COLUNA 6
tmp(56) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(57) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(58) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(59) := "11" & x"4" & '0' & x"0F";	-- LDI 15, R3	#O
tmp(60) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(61) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(62) := "11" & x"4" & '0' & x"07";	-- LDI 7, R3	#COLUNA 7
tmp(63) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(64) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(65) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(66) := "11" & x"4" & '0' & x"07";	-- LDI 7, R3	#G
tmp(67) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(68) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(69) := "11" & x"4" & '0' & x"08";	-- LDI 8, R3	#COLUNA 8
tmp(70) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(71) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(72) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(73) := "11" & x"4" & '0' & x"09";	-- LDI 9, R3	#I
tmp(74) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(75) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(76) := "11" & x"4" & '0' & x"09";	-- LDI 9, R3	#COLUNA 9
tmp(77) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(78) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(79) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(80) := "11" & x"4" & '0' & x"0F";	-- LDI 15, R3	#O
tmp(81) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(82) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(83) := "11" & x"4" & '0' & x"0B";	-- LDI 11, R3	#COLUNA 11
tmp(84) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(85) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(86) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(87) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#B
tmp(88) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(89) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(90) := "11" & x"4" & '0' & x"0C";	-- LDI 12, R3	#COLUNA 12
tmp(91) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(92) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(93) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(94) := "11" & x"4" & '0' & x"01";	-- LDI 1, R3	#A
tmp(95) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(96) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(97) := "11" & x"4" & '0' & x"0D";	-- LDI 13, R3	#COLUNA 13
tmp(98) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(99) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(100) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(101) := "11" & x"4" & '0' & x"03";	-- LDI 3, R3	#C
tmp(102) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(103) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(104) := "11" & x"4" & '0' & x"0E";	-- LDI 14, R3	#COLUNA 14
tmp(105) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(106) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(107) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(108) := "11" & x"4" & '0' & x"01";	-- LDI 1, R3	#A
tmp(109) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(110) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(111) := "11" & x"4" & '0' & x"0F";	-- LDI 15, R3	#COLUNA 15
tmp(112) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(113) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(114) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(115) := "11" & x"4" & '0' & x"0E";	-- LDI 14, R3	#N
tmp(116) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(117) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(118) := "11" & x"4" & '0' & x"10";	-- LDI 16, R3	#COLUNA 16
tmp(119) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(120) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(121) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(122) := "11" & x"4" & '0' & x"01";	-- LDI 1, R3	#A
tmp(123) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(124) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(125) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(126) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(127) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(128) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(129) := "00" & x"1" & '1' & x"60";	-- LDA 352, R0	#Carrega o acumulador com a leitura do botão KEY0
tmp(130) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(131) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(132) := "00" & x"7" & '0' & x"87";	-- JEQ NAO_CLICOU0	#Desvia se igual a 0 (botão não foi pressionado)
tmp(133) := "00" & x"9" & '0' & x"9F";	-- JSR INCREMENTO	#O botão foi pressionado, chama a sub-rotina de incremento
tmp(134) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de incremento
tmp(135) := "00" & x"9" & '0' & x"D8";	-- JSR SALVA_DISP	#Escreve o valor das váriaveis de contagem nos displays
tmp(136) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de salvar nos displays
tmp(137) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(138) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(139) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(140) := "00" & x"7" & '0' & x"8F";	-- JEQ NAO_CLICOU1	#Desvia se igual a 0 (botão não foi pressionado)
tmp(141) := "00" & x"9" & '1' & x"12";	-- JSR DEFINE_LIM	#O botão foi pressionado, chama a sub-rotina de incremento
tmp(142) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de definir limite
tmp(143) := "00" & x"9" & '0' & x"F6";	-- JSR VERIFICA_LIM
tmp(144) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de verificar limite
tmp(145) := "00" & x"1" & '1' & x"62";	-- LDA 354, R0	#Carrega o acumulador com a leitura do botão KEY2
tmp(146) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(147) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(148) := "00" & x"7" & '0' & x"97";	-- JEQ NAO_CLICOU2	#Desvia se igual a 0 (botão não foi pressionado)
tmp(149) := "00" & x"9" & '1' & x"47";	-- JSR DECREMENTO	#O botão foi pressionado, chama a sub-rotina de incremento
tmp(150) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de incremento
tmp(151) := "00" & x"1" & '1' & x"64";	-- LDA 356, R0	#Carrega o acumulador com a leitura do botão FPGA_RESET
tmp(152) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(153) := "00" & x"D" & '0' & x"01";	-- CEQi 1, R0	#Compara com constante 1
tmp(154) := "00" & x"7" & '0' & x"9C";	-- JEQ REINICIO	#Desvia se igual a 1 (botão não foi pressionado)
tmp(155) := "00" & x"9" & '0' & x"E5";	-- JSR RESET	#O botão foi pressionado, chama a sub-rotina de reset
tmp(156) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de reset
tmp(157) := "00" & x"6" & '0' & x"80";	-- JMP INICIO	#Fecha o laço principal, faz uma nova leitura de KEY0
tmp(158) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(159) := "00" & x"5" & '1' & x"FF";	-- STA 511, R0	#Limpa a leitura do botão
tmp(160) := "00" & x"1" & '0' & x"09";	-- LDA 9, R0	#Carrega o valor de MEM[9] (flag inibir contagem)
tmp(161) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara o valor com constante 0
tmp(162) := "00" & x"7" & '0' & x"A4";	-- JEQ INCREMENTAR
tmp(163) := "00" & x"A" & '0' & x"00";	-- RET
tmp(164) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	#Carrega o valor de MEM[0] (contador)
tmp(165) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(166) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(167) := "00" & x"7" & '0' & x"AA";	-- JEQ VAIUM_D	#Realiza o carry out caso valor igual a 10
tmp(168) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Salva o incremento em MEM[0] (contador)
tmp(169) := "00" & x"A" & '0' & x"00";	-- RET	#Retorna da sub-rotina
tmp(170) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(171) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador em MEM[0] (unidades)
tmp(172) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	#Carrega valor de MEM[1] no acumulador (dezenas)
tmp(173) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(174) := "00" & x"D" & '0' & x"06";	-- CEQi 6, R0	#Compara o valor com constante 10
tmp(175) := "00" & x"7" & '0' & x"B2";	-- JEQ VAIUM_C	#Realiza o carry out caso valor igual a 10
tmp(176) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Salva o incremento em MEM[1] (dezenas)
tmp(177) := "00" & x"A" & '0' & x"00";	-- RET
tmp(178) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(179) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador em MEM[1] (dezenas)
tmp(180) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	#Carrega valor de MEM[2] no acumulador (centenas)
tmp(181) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(182) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(183) := "00" & x"7" & '0' & x"BA";	-- JEQ VAIUM_M	#Realiza o carry out caso valor igual a 10
tmp(184) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Salva o incremento em MEM[2] (centenas)
tmp(185) := "00" & x"A" & '0' & x"00";	-- RET
tmp(186) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(187) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador em MEM[2] (centenas)
tmp(188) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	#Carrega valor de MEM[6] no acumulador (milhares)
tmp(189) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(190) := "00" & x"D" & '0' & x"06";	-- CEQi 6, R0	#Compara o valor com constante 10
tmp(191) := "00" & x"7" & '0' & x"C2";	-- JEQ VAIUM_DM	#Realiza o carry out caso valor igual a 10
tmp(192) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Salva o incremento em MEM[6] (milhares)
tmp(193) := "00" & x"A" & '0' & x"00";	-- RET
tmp(194) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(195) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador em MEM[6] (milhares)
tmp(196) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	#Carrega valor de MEM[7] no acumulador (dezenas de milhares)
tmp(197) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(198) := "01" & x"1" & '0' & x"08";	-- LDA 8, R1	#Carrega valor de MEM[8] no acumulador (centenas de milhares)
tmp(199) := "01" & x"D" & '0' & x"02";	-- CEQi 2, R1	#Compara o valor com constante 2
tmp(200) := "00" & x"7" & '0' & x"CC";	-- JEQ COMPARA4	#Pula para o fim da rotina
tmp(201) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(202) := "00" & x"7" & '0' & x"D0";	-- JEQ VAIUM_CM	#Realiza o carry out caso valor igual a 10
tmp(203) := "00" & x"6" & '0' & x"CE";	-- JMP END_DM
tmp(204) := "00" & x"D" & '0' & x"04";	-- CEQi 4, R0	#Compara o valor com constante 4
tmp(205) := "00" & x"7" & '0' & x"D0";	-- JEQ VAIUM_CM	#Realiza o carry out caso valor igual a 4
tmp(206) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Salva o incremento em MEM[7] (dezenas de milhares)
tmp(207) := "00" & x"A" & '0' & x"00";	-- RET
tmp(208) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(209) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador em MEM[7] (dezenas milhares)
tmp(210) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega valor de MEM[8] no acumulador (centenas de milhares)
tmp(211) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(212) := "00" & x"D" & '0' & x"03";	-- CEQi 3, R0	#Compara o valor com constante 3
tmp(213) := "00" & x"7" & '1' & x"79";	-- JEQ ZERA_HEX	#Zera se chegar ao final
tmp(214) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Salva o incremento em MEM[8] (centena de milhares)
tmp(215) := "00" & x"A" & '0' & x"00";	-- RET
tmp(216) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	#Carrega o valor de MEM[0] (unidades)
tmp(217) := "00" & x"5" & '1' & x"20";	-- STA 288, R0	#Armazena valor do acumulador de unidades no HEX0
tmp(218) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	#Carrega o valor de MEM[1] (dezenas)
tmp(219) := "00" & x"5" & '1' & x"21";	-- STA 289, R0	#Armazena valor do acumulador de dezenas no HEX1
tmp(220) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	#Carrega o valor de MEM[2] (centenas)
tmp(221) := "00" & x"5" & '1' & x"22";	-- STA 290, R0	#Armazena valor do acumulador de centenas no HEX2
tmp(222) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	#Carrega o valor de MEM[6] (milhares)
tmp(223) := "00" & x"5" & '1' & x"23";	-- STA 291, R0	#Armazena valor do acumulador de unidades no HEX3
tmp(224) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	#Carrega o valor de MEM[7] (dezenas de milhares)
tmp(225) := "00" & x"5" & '1' & x"24";	-- STA 292, R0	#Armazena valor do acumulador de dezenas no HEX4
tmp(226) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega o valor de MEM[8] (centenas de milhares)
tmp(227) := "00" & x"5" & '1' & x"25";	-- STA 293, R0	#Armazena valor do acumulador de centenas no HEX5
tmp(228) := "00" & x"A" & '0' & x"00";	-- RET
tmp(229) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(230) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador na MEM[0] (unidades)
tmp(231) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador na MEM[1] (dezenas)
tmp(232) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador na MEM[2] (centenas)
tmp(233) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador na MEM[6] (milhar)
tmp(234) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador na MEM[7] (dezena de milhar)
tmp(235) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do acumulador na MEM[8] (centena de milhar)
tmp(236) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador na MEM[9] (flag inibir contagem)
tmp(237) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(238) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega o acumulador com o valor 9
tmp(239) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do acumulador em MEM[10] (inibir unidade)
tmp(240) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do acumulador em MEM[11] (inibir dezena)
tmp(241) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do acumulador em MEM[12] (inibir centena)
tmp(242) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do acumulador em MEM[13] (inibir milhar)
tmp(243) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do acumulador em MEM[14] (inibir dezena de milhar)
tmp(244) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do acumulador em MEM[15] (inibir centena de milhar)
tmp(245) := "00" & x"A" & '0' & x"00";	-- RET
tmp(246) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	#Carrega o valor de MEM[0] (unidades)
tmp(247) := "00" & x"8" & '0' & x"0A";	-- CEQ 10, R0	#Compara o valor de MEM[10] (inibir unidade)
tmp(248) := "00" & x"7" & '0' & x"FA";	-- JEQ NEXT_LIM1
tmp(249) := "00" & x"A" & '0' & x"00";	-- RET
tmp(250) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	#Carrega o valor de MEM[1] (dezenas)
tmp(251) := "00" & x"8" & '0' & x"0B";	-- CEQ 11, R0	#Compara o valor de MEM[11] (inibir dezenas)
tmp(252) := "00" & x"7" & '0' & x"FE";	-- JEQ NEXT_LIM2
tmp(253) := "00" & x"A" & '0' & x"00";	-- RET
tmp(254) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	#Carrega o valor de MEM[2] (centenas)
tmp(255) := "00" & x"8" & '0' & x"0C";	-- CEQ 12, R0	#Compara o valor de MEM[12] (inibir centenas)
tmp(256) := "00" & x"7" & '1' & x"02";	-- JEQ NEXT_LIM3
tmp(257) := "00" & x"A" & '0' & x"00";	-- RET
tmp(258) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	#Carrega o valor de MEM[6] (milhar)
tmp(259) := "00" & x"8" & '0' & x"0D";	-- CEQ 13, R0	#Compara o valor de MEM[13] (inibir milhar)
tmp(260) := "00" & x"7" & '1' & x"06";	-- JEQ NEXT_LIM4
tmp(261) := "00" & x"A" & '0' & x"00";	-- RET
tmp(262) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	#Carrega o valor de MEM[7] (dezena de milhar)
tmp(263) := "00" & x"8" & '0' & x"0E";	-- CEQ 14, R0	#Compara o valor de MEM[10] (inibir dezena de milhar)
tmp(264) := "00" & x"7" & '1' & x"0A";	-- JEQ NEXT_LIM5
tmp(265) := "00" & x"A" & '0' & x"00";	-- RET
tmp(266) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega o valor de MEM[8] (centena de milhar)
tmp(267) := "00" & x"8" & '0' & x"0F";	-- CEQ 15, R0	#Compara o valor de MEM[10] (inibir centena de milhar)
tmp(268) := "00" & x"7" & '1' & x"0E";	-- JEQ TODOS_IGUAL
tmp(269) := "00" & x"A" & '0' & x"00";	-- RET
tmp(270) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o acumulador com o valor 1
tmp(271) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador em MEM[9] (flag inibir contagem)
tmp(272) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(273) := "00" & x"A" & '0' & x"00";	-- RET
tmp(274) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(275) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(276) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do acumulador em MEM[10] (inibir unidade)
tmp(277) := "00" & x"4" & '0' & x"04";	-- LDI 4, R0	#Carrega o acumulador com o valor 4
tmp(278) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(279) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(280) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(281) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(282) := "00" & x"7" & '1' & x"17";	-- JEQ AGUARDA_D	#Desvia se igual a 0 (botão não foi pressionado)
tmp(283) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(284) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(285) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do acumulador em MEM[11] (inibir dezena)
tmp(286) := "00" & x"4" & '0' & x"10";	-- LDI 16, R0	#Carrega o acumulador com o valor 16
tmp(287) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(288) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(289) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(290) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(291) := "00" & x"7" & '1' & x"20";	-- JEQ AGUARDA_C	#Desvia se igual a 0 (botão não foi pressionado)
tmp(292) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(293) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(294) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do acumulador em MEM[12] (inibir centena)
tmp(295) := "00" & x"4" & '0' & x"20";	-- LDI 32, R0	#Carrega o acumulador com o valor 32
tmp(296) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(297) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(298) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(299) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(300) := "00" & x"7" & '1' & x"29";	-- JEQ AGUARDA_M	#Desvia se igual a 0 (botão não foi pressionado)
tmp(301) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(302) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(303) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do acumulador em MEM[13] (inibir milhar)
tmp(304) := "00" & x"4" & '0' & x"80";	-- LDI 128, R0	#Carrega o acumulador com o valor 128
tmp(305) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(306) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(307) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(308) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(309) := "00" & x"7" & '1' & x"32";	-- JEQ AGUARDA_DM	#Desvia se igual a 0 (botão não foi pressionado)
tmp(310) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(311) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(312) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do acumulador em MEM[13] (inibir dezena de milhar)
tmp(313) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(314) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(315) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o acumulador com o valor 1
tmp(316) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do acumulador no LDR9
tmp(317) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(318) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(319) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(320) := "00" & x"7" & '1' & x"3D";	-- JEQ AGUARDA_CM	#Desvia se igual a 0 (botão não foi pressionado)
tmp(321) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(322) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(323) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do acumulador em MEM[15] (inibir centena de milhar)
tmp(324) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(325) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do acumulador no LDR9
tmp(326) := "00" & x"A" & '0' & x"00";	-- RET
tmp(327) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega 0 para o acumulador
tmp(328) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(329) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador na MEM[9] (flag inibir contagem)
tmp(330) := "00" & x"5" & '1' & x"FD";	-- STA 509, R0	#Limpa a leitura do botão KEY2
tmp(331) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	# Carrega MEM[0] (unidades) no acumulador
tmp(332) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[0] == 0
tmp(333) := "00" & x"7" & '1' & x"51";	-- JEQ VEMUM_D	# Se MEM[0] == 0, realiza o "empréstimo"
tmp(334) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[0]
tmp(335) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	# Armazena o novo valor de MEM[0]
tmp(336) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(337) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(338) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	# Define MEM[0] para 9
tmp(339) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	# Carrega MEM[1] (dezenas) no acumulador
tmp(340) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[1] == 0
tmp(341) := "00" & x"7" & '1' & x"59";	-- JEQ VEMUM_C	# Se MEM[1] == 0, realiza o próximo "empréstimo"
tmp(342) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[1]
tmp(343) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	# Armazena o novo valor de MEM[1]
tmp(344) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(345) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(346) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	# Define MEM[1] para 9
tmp(347) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	# Carrega MEM[2] (centenas) no acumulador
tmp(348) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[2] == 0
tmp(349) := "00" & x"7" & '1' & x"61";	-- JEQ VEMUM_M	# Se MEM[2] == 0, realiza o próximo "empréstimo"
tmp(350) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[2]
tmp(351) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	# Armazena o novo valor de MEM[2]
tmp(352) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(353) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(354) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	# Define MEM[2] para 9
tmp(355) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	# Carrega MEM[3] (milhares) no acumulador
tmp(356) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[3] == 0
tmp(357) := "00" & x"7" & '1' & x"69";	-- JEQ VEMUM_DM	# Se MEM[3] == 0, realiza o próximo "empréstimo"
tmp(358) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[3]
tmp(359) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	# Armazena o novo valor de MEM[3]
tmp(360) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(361) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(362) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	# Define MEM[3] para 9
tmp(363) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	# Carrega MEM[4] (dezenas de milhares) no acumulador
tmp(364) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[4] == 0
tmp(365) := "00" & x"7" & '1' & x"71";	-- JEQ VEMUM_CM	# Se MEM[4] == 0, realiza o próximo "empréstimo"
tmp(366) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[4]
tmp(367) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	# Armazena o novo valor de MEM[4]
tmp(368) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(369) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(370) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	# Define MEM[4] para 9
tmp(371) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	# Carrega MEM[5] (centenas de milhares) no acumulador
tmp(372) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[5] == 0
tmp(373) := "00" & x"7" & '1' & x"79";	-- JEQ ZERA_HEX	# Zera se for menos que 0
tmp(374) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[5]
tmp(375) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	# Armazena o novo valor de MEM[5]
tmp(376) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(377) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(378) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador na MEM[0] (unidades)
tmp(379) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador na MEM[1] (dezenas)
tmp(380) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador na MEM[2] (centenas)
tmp(381) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador na MEM[6] (milhar)
tmp(382) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador na MEM[7] (dezena de milhar)
tmp(383) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do acumulador na MEM[8] (centena de milhar)
tmp(384) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador na MEM[9] (flag inibir contagem)
tmp(385) := "00" & x"A" & '0' & x"00";	-- RET


        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;