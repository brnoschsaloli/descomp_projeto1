library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Operacao_ULA_2bits, habLeituraMEM, habEscritaMEM 
      -- Inicializa os endereços:
tmp(0) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(1) := "00" & x"5" & '1' & x"20";	-- STA 288, R0	#Armazena o valor do acumulador em HEX0
tmp(2) := "00" & x"5" & '1' & x"21";	-- STA 289, R0	#Armazena o valor do acumulador em HEX1
tmp(3) := "00" & x"5" & '1' & x"22";	-- STA 290, R0	#Armazena o valor do acumulador em HEX2
tmp(4) := "00" & x"5" & '1' & x"23";	-- STA 291, R0	#Armazena o valor do acumulador em HEX3
tmp(5) := "00" & x"5" & '1' & x"24";	-- STA 292, R0	#Armazena o valor do acumulador em HEX4
tmp(6) := "00" & x"5" & '1' & x"25";	-- STA 293, R0	#Armazena o valor do acumulador em HEX5
tmp(7) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(8) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(9) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(10) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(11) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do acumulador no LDR9
tmp(12) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(13) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(14) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador em MEM[0] (unidades)
tmp(15) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador em MEM[1] (dezenas)
tmp(16) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador em MEM[2] (centenas)
tmp(17) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador em MEM[6] (milhares)
tmp(18) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador em MEM[7] (dezenas de milhares)
tmp(19) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do acumulador em MEM[8] (centenas de milhares)
tmp(20) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador em MEM[9] (flag inibir contagem)
tmp(21) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega o acumulador com o valor 9
tmp(22) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do acumulador em MEM[10] (inibir unidade)
tmp(23) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do acumulador em MEM[11] (inibir dezena)
tmp(24) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do acumulador em MEM[12] (inibir centena)
tmp(25) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do acumulador em MEM[13] (inibir milhar)
tmp(26) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do acumulador em MEM[14] (inibir dezena de milhar)
tmp(27) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do acumulador em MEM[15] (inibir centena de milhar)
tmp(28) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(29) := "00" & x"5" & '1' & x"FF";	-- STA 511, R0	#Limpa a leitura do botão zero
tmp(30) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(31) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(32) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(33) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(34) := "11" & x"4" & '0' & x"03";	-- LDI 3, R3	#COLUNA 3
tmp(35) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(36) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(37) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(38) := "11" & x"4" & '0' & x"10";	-- LDI 16, R3	#P
tmp(39) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(40) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(41) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#COLUNA 4
tmp(42) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(43) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(44) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(45) := "11" & x"4" & '0' & x"01";	-- LDI 1, R3	#A
tmp(46) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(47) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(48) := "11" & x"4" & '0' & x"05";	-- LDI 5, R3	#COLUNA 5
tmp(49) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(50) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(51) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(52) := "11" & x"4" & '0' & x"15";	-- LDI 21, R3	#U
tmp(53) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(54) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(55) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#COLUNA 6
tmp(56) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(57) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(58) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(59) := "11" & x"4" & '0' & x"0C";	-- LDI 12, R3	#L
tmp(60) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(61) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(62) := "11" & x"4" & '0' & x"07";	-- LDI 7, R3	#COLUNA 7
tmp(63) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(64) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(65) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(66) := "11" & x"4" & '0' & x"01";	-- LDI 1, R3	#A
tmp(67) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(68) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(69) := "11" & x"4" & '0' & x"08";	-- LDI 8, R3	#COLUNA 8
tmp(70) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(71) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(72) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(73) := "11" & x"4" & '0' & x"0F";	-- LDI 15, R3	#O
tmp(74) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(75) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(76) := "11" & x"4" & '0' & x"0A";	-- LDI 10, R3	#COLUNA 10
tmp(77) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(78) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(79) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(80) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#B
tmp(81) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(82) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(83) := "11" & x"4" & '0' & x"0B";	-- LDI 11, R3	#COLUNA 11
tmp(84) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(85) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(86) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(87) := "11" & x"4" & '0' & x"0F";	-- LDI 15, R3	#O
tmp(88) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(89) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(90) := "11" & x"4" & '0' & x"0C";	-- LDI 12, R3	#COLUNA 12
tmp(91) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(92) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(93) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(94) := "11" & x"4" & '0' & x"0E";	-- LDI 14, R3	#N
tmp(95) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(96) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(97) := "11" & x"4" & '0' & x"0D";	-- LDI 13, R3	#COLUNA 13
tmp(98) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(99) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(100) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(101) := "11" & x"4" & '0' & x"09";	-- LDI 9, R3	#I
tmp(102) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(103) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(104) := "11" & x"4" & '0' & x"0E";	-- LDI 14, R3	#COLUNA 14
tmp(105) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(106) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(107) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(108) := "11" & x"4" & '0' & x"14";	-- LDI 20, R3	#T
tmp(109) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(110) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(111) := "11" & x"4" & '0' & x"0F";	-- LDI 15, R3	#COLUNA 15
tmp(112) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(113) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(114) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(115) := "11" & x"4" & '0' & x"01";	-- LDI 1, R3	#A
tmp(116) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(117) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(118) := "11" & x"4" & '0' & x"10";	-- LDI 16, R3	#COLUNA 16
tmp(119) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(120) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(121) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(122) := "11" & x"4" & '0' & x"0F";	-- LDI 15, R3	#O
tmp(123) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(124) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(125) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(126) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(127) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(128) := "11" & x"4" & '0' & x"08";	-- LDI 8, R3	#COLUNA 8
tmp(129) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(130) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(131) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(132) := "11" & x"4" & '0' & x"3A";	-- LDI 58, R3	#dois pontos
tmp(133) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(134) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(135) := "11" & x"4" & '0' & x"0B";	-- LDI 11, R3	#COLUNA 11
tmp(136) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(137) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(138) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(139) := "11" & x"4" & '0' & x"3A";	-- LDI 58, R3	#dois pontos
tmp(140) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(141) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(142) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(143) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(144) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(145) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(146) := "00" & x"1" & '1' & x"60";	-- LDA 352, R0	#Carrega o acumulador com a leitura do botão KEY0
tmp(147) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(148) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(149) := "00" & x"7" & '0' & x"98";	-- JEQ NAO_CLICOU0	#Desvia se igual a 0 (botão não foi pressionado)
tmp(150) := "00" & x"9" & '0' & x"B0";	-- JSR INCREMENTO	#O botão foi pressionado, chama a sub-rotina de incremento
tmp(151) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de incremento
tmp(152) := "00" & x"9" & '0' & x"E9";	-- JSR SALVA_DISP	#Escreve o valor das váriaveis de contagem nos displays
tmp(153) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de salvar nos displays
tmp(154) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(155) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(156) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(157) := "00" & x"7" & '0' & x"A0";	-- JEQ NAO_CLICOU1	#Desvia se igual a 0 (botão não foi pressionado)
tmp(158) := "00" & x"9" & '1' & x"53";	-- JSR DEFINE_LIM	#O botão foi pressionado, chama a sub-rotina de incremento
tmp(159) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de definir limite
tmp(160) := "00" & x"9" & '1' & x"37";	-- JSR VERIFICA_LIM
tmp(161) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de verificar limite
tmp(162) := "00" & x"1" & '1' & x"62";	-- LDA 354, R0	#Carrega o acumulador com a leitura do botão KEY2
tmp(163) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(164) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(165) := "00" & x"7" & '0' & x"A8";	-- JEQ NAO_CLICOU2	#Desvia se igual a 0 (botão não foi pressionado)
tmp(166) := "00" & x"9" & '1' & x"88";	-- JSR DECREMENTO	#O botão foi pressionado, chama a sub-rotina de incremento
tmp(167) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de incremento
tmp(168) := "00" & x"1" & '1' & x"64";	-- LDA 356, R0	#Carrega o acumulador com a leitura do botão FPGA_RESET
tmp(169) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(170) := "00" & x"D" & '0' & x"01";	-- CEQi 1, R0	#Compara com constante 1
tmp(171) := "00" & x"7" & '0' & x"AD";	-- JEQ REINICIO	#Desvia se igual a 1 (botão não foi pressionado)
tmp(172) := "00" & x"9" & '1' & x"26";	-- JSR RESET	#O botão foi pressionado, chama a sub-rotina de reset
tmp(173) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de reset
tmp(174) := "00" & x"6" & '0' & x"91";	-- JMP INICIO	#Fecha o laço principal, faz uma nova leitura de KEY0
tmp(175) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(176) := "00" & x"5" & '1' & x"FF";	-- STA 511, R0	#Limpa a leitura do botão
tmp(177) := "00" & x"1" & '0' & x"09";	-- LDA 9, R0	#Carrega o valor de MEM[9] (flag inibir contagem)
tmp(178) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara o valor com constante 0
tmp(179) := "00" & x"7" & '0' & x"B5";	-- JEQ INCREMENTAR
tmp(180) := "00" & x"A" & '0' & x"00";	-- RET
tmp(181) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	#Carrega o valor de MEM[0] (contador)
tmp(182) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(183) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(184) := "00" & x"7" & '0' & x"BB";	-- JEQ VAIUM_D	#Realiza o carry out caso valor igual a 10
tmp(185) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Salva o incremento em MEM[0] (contador)
tmp(186) := "00" & x"A" & '0' & x"00";	-- RET	#Retorna da sub-rotina
tmp(187) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(188) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador em MEM[0] (unidades)
tmp(189) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	#Carrega valor de MEM[1] no acumulador (dezenas)
tmp(190) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(191) := "00" & x"D" & '0' & x"06";	-- CEQi 6, R0	#Compara o valor com constante 10
tmp(192) := "00" & x"7" & '0' & x"C3";	-- JEQ VAIUM_C	#Realiza o carry out caso valor igual a 10
tmp(193) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Salva o incremento em MEM[1] (dezenas)
tmp(194) := "00" & x"A" & '0' & x"00";	-- RET
tmp(195) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(196) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador em MEM[1] (dezenas)
tmp(197) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	#Carrega valor de MEM[2] no acumulador (centenas)
tmp(198) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(199) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(200) := "00" & x"7" & '0' & x"CB";	-- JEQ VAIUM_M	#Realiza o carry out caso valor igual a 10
tmp(201) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Salva o incremento em MEM[2] (centenas)
tmp(202) := "00" & x"A" & '0' & x"00";	-- RET
tmp(203) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(204) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador em MEM[2] (centenas)
tmp(205) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	#Carrega valor de MEM[6] no acumulador (milhares)
tmp(206) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(207) := "00" & x"D" & '0' & x"06";	-- CEQi 6, R0	#Compara o valor com constante 10
tmp(208) := "00" & x"7" & '0' & x"D3";	-- JEQ VAIUM_DM	#Realiza o carry out caso valor igual a 10
tmp(209) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Salva o incremento em MEM[6] (milhares)
tmp(210) := "00" & x"A" & '0' & x"00";	-- RET
tmp(211) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(212) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador em MEM[6] (milhares)
tmp(213) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	#Carrega valor de MEM[7] no acumulador (dezenas de milhares)
tmp(214) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(215) := "01" & x"1" & '0' & x"08";	-- LDA 8, R1	#Carrega valor de MEM[8] no acumulador (centenas de milhares)
tmp(216) := "01" & x"D" & '0' & x"02";	-- CEQi 2, R1	#Compara o valor com constante 2
tmp(217) := "00" & x"7" & '0' & x"DD";	-- JEQ COMPARA4	#Pula para o fim da rotina
tmp(218) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(219) := "00" & x"7" & '0' & x"E1";	-- JEQ VAIUM_CM	#Realiza o carry out caso valor igual a 10
tmp(220) := "00" & x"6" & '0' & x"DF";	-- JMP END_DM
tmp(221) := "00" & x"D" & '0' & x"04";	-- CEQi 4, R0	#Compara o valor com constante 4
tmp(222) := "00" & x"7" & '0' & x"E1";	-- JEQ VAIUM_CM	#Realiza o carry out caso valor igual a 4
tmp(223) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Salva o incremento em MEM[7] (dezenas de milhares)
tmp(224) := "00" & x"A" & '0' & x"00";	-- RET
tmp(225) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(226) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador em MEM[7] (dezenas milhares)
tmp(227) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega valor de MEM[8] no acumulador (centenas de milhares)
tmp(228) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(229) := "00" & x"D" & '0' & x"03";	-- CEQi 3, R0	#Compara o valor com constante 3
tmp(230) := "00" & x"7" & '1' & x"BA";	-- JEQ ZERA_HEX	#Zera se chegar ao final
tmp(231) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Salva o incremento em MEM[8] (centena de milhares)
tmp(232) := "00" & x"A" & '0' & x"00";	-- RET
tmp(233) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(234) := "11" & x"4" & '0' & x"0D";	-- LDI 13, R3	#COLUNA 13
tmp(235) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(236) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(237) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(238) := "11" & x"1" & '0' & x"00";	-- LDA 0, R3	#Carrega o valor de MEM[0] (unidades)
tmp(239) := "11" & x"5" & '1' & x"20";	-- STA 288, R3	#Armazena valor do acumulador de unidades no HEX0
tmp(240) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(241) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(242) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(243) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(244) := "11" & x"4" & '0' & x"0C";	-- LDI 12, R3	#COLUNA 12
tmp(245) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(246) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(247) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(248) := "11" & x"1" & '0' & x"01";	-- LDA 1, R3	#Carrega o valor de MEM[1] (dezenas)
tmp(249) := "11" & x"5" & '1' & x"21";	-- STA 289, R3	#Armazena valor do acumulador de dezenas no HEX1
tmp(250) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(251) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(252) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(253) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(254) := "11" & x"4" & '0' & x"0A";	-- LDI 10, R3	#COLUNA 10
tmp(255) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(256) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(257) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(258) := "11" & x"1" & '0' & x"02";	-- LDA 2, R3	#Carrega o valor de MEM[2] (centenas)
tmp(259) := "11" & x"5" & '1' & x"22";	-- STA 290, R3	#Armazena valor do acumulador de centenas no HEX2
tmp(260) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(261) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(262) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(263) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(264) := "11" & x"4" & '0' & x"09";	-- LDI 9, R3	#COLUNA 9
tmp(265) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(266) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(267) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(268) := "11" & x"1" & '0' & x"06";	-- LDA 6, R3	#Carrega o valor de MEM[6] (milhares)
tmp(269) := "11" & x"5" & '1' & x"23";	-- STA 291, R3	#Armazena valor do acumulador de unidades no HEX3
tmp(270) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(271) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(272) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(273) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(274) := "11" & x"4" & '0' & x"07";	-- LDI 7, R3	#COLUNA 7
tmp(275) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(276) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(277) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(278) := "11" & x"1" & '0' & x"07";	-- LDA 7, R3	#Carrega o valor de MEM[7] (dezenas de milhares)
tmp(279) := "11" & x"5" & '1' & x"24";	-- STA 292, R3	#Armazena valor do acumulador de dezenas no HEX4
tmp(280) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(281) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(282) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(283) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(284) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#COLUNA 6
tmp(285) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(286) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(287) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(288) := "11" & x"1" & '0' & x"08";	-- LDA 8, R3	#Carrega o valor de MEM[8] (centenas de milhares)
tmp(289) := "11" & x"5" & '1' & x"25";	-- STA 293, R3	#Armazena valor do acumulador de centenas no HEX5
tmp(290) := "11" & x"E" & '0' & x"30";	-- ADDi 48, R3	#ACERTA COM O VALOR NO DO NUMERO NO .MIF
tmp(291) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(292) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(293) := "00" & x"A" & '0' & x"00";	-- RET
tmp(294) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(295) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador na MEM[0] (unidades)
tmp(296) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador na MEM[1] (dezenas)
tmp(297) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador na MEM[2] (centenas)
tmp(298) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador na MEM[6] (milhar)
tmp(299) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador na MEM[7] (dezena de milhar)
tmp(300) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do acumulador na MEM[8] (centena de milhar)
tmp(301) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador na MEM[9] (flag inibir contagem)
tmp(302) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(303) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega o acumulador com o valor 9
tmp(304) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do acumulador em MEM[10] (inibir unidade)
tmp(305) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do acumulador em MEM[11] (inibir dezena)
tmp(306) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do acumulador em MEM[12] (inibir centena)
tmp(307) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do acumulador em MEM[13] (inibir milhar)
tmp(308) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do acumulador em MEM[14] (inibir dezena de milhar)
tmp(309) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do acumulador em MEM[15] (inibir centena de milhar)
tmp(310) := "00" & x"A" & '0' & x"00";	-- RET
tmp(311) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	#Carrega o valor de MEM[0] (unidades)
tmp(312) := "00" & x"8" & '0' & x"0A";	-- CEQ 10, R0	#Compara o valor de MEM[10] (inibir unidade)
tmp(313) := "00" & x"7" & '1' & x"3B";	-- JEQ NEXT_LIM1
tmp(314) := "00" & x"A" & '0' & x"00";	-- RET
tmp(315) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	#Carrega o valor de MEM[1] (dezenas)
tmp(316) := "00" & x"8" & '0' & x"0B";	-- CEQ 11, R0	#Compara o valor de MEM[11] (inibir dezenas)
tmp(317) := "00" & x"7" & '1' & x"3F";	-- JEQ NEXT_LIM2
tmp(318) := "00" & x"A" & '0' & x"00";	-- RET
tmp(319) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	#Carrega o valor de MEM[2] (centenas)
tmp(320) := "00" & x"8" & '0' & x"0C";	-- CEQ 12, R0	#Compara o valor de MEM[12] (inibir centenas)
tmp(321) := "00" & x"7" & '1' & x"43";	-- JEQ NEXT_LIM3
tmp(322) := "00" & x"A" & '0' & x"00";	-- RET
tmp(323) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	#Carrega o valor de MEM[6] (milhar)
tmp(324) := "00" & x"8" & '0' & x"0D";	-- CEQ 13, R0	#Compara o valor de MEM[13] (inibir milhar)
tmp(325) := "00" & x"7" & '1' & x"47";	-- JEQ NEXT_LIM4
tmp(326) := "00" & x"A" & '0' & x"00";	-- RET
tmp(327) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	#Carrega o valor de MEM[7] (dezena de milhar)
tmp(328) := "00" & x"8" & '0' & x"0E";	-- CEQ 14, R0	#Compara o valor de MEM[10] (inibir dezena de milhar)
tmp(329) := "00" & x"7" & '1' & x"4B";	-- JEQ NEXT_LIM5
tmp(330) := "00" & x"A" & '0' & x"00";	-- RET
tmp(331) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega o valor de MEM[8] (centena de milhar)
tmp(332) := "00" & x"8" & '0' & x"0F";	-- CEQ 15, R0	#Compara o valor de MEM[10] (inibir centena de milhar)
tmp(333) := "00" & x"7" & '1' & x"4F";	-- JEQ TODOS_IGUAL
tmp(334) := "00" & x"A" & '0' & x"00";	-- RET
tmp(335) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o acumulador com o valor 1
tmp(336) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador em MEM[9] (flag inibir contagem)
tmp(337) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(338) := "00" & x"A" & '0' & x"00";	-- RET
tmp(339) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(340) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(341) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do acumulador em MEM[10] (inibir unidade)
tmp(342) := "00" & x"4" & '0' & x"04";	-- LDI 4, R0	#Carrega o acumulador com o valor 4
tmp(343) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(344) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(345) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(346) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(347) := "00" & x"7" & '1' & x"58";	-- JEQ AGUARDA_D	#Desvia se igual a 0 (botão não foi pressionado)
tmp(348) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(349) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(350) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do acumulador em MEM[11] (inibir dezena)
tmp(351) := "00" & x"4" & '0' & x"10";	-- LDI 16, R0	#Carrega o acumulador com o valor 16
tmp(352) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(353) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(354) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(355) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(356) := "00" & x"7" & '1' & x"61";	-- JEQ AGUARDA_C	#Desvia se igual a 0 (botão não foi pressionado)
tmp(357) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(358) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(359) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do acumulador em MEM[12] (inibir centena)
tmp(360) := "00" & x"4" & '0' & x"20";	-- LDI 32, R0	#Carrega o acumulador com o valor 32
tmp(361) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(362) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(363) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(364) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(365) := "00" & x"7" & '1' & x"6A";	-- JEQ AGUARDA_M	#Desvia se igual a 0 (botão não foi pressionado)
tmp(366) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(367) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(368) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do acumulador em MEM[13] (inibir milhar)
tmp(369) := "00" & x"4" & '0' & x"80";	-- LDI 128, R0	#Carrega o acumulador com o valor 128
tmp(370) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(371) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(372) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(373) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(374) := "00" & x"7" & '1' & x"73";	-- JEQ AGUARDA_DM	#Desvia se igual a 0 (botão não foi pressionado)
tmp(375) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(376) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(377) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do acumulador em MEM[13] (inibir dezena de milhar)
tmp(378) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(379) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(380) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o acumulador com o valor 1
tmp(381) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do acumulador no LDR9
tmp(382) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(383) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(384) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(385) := "00" & x"7" & '1' & x"7E";	-- JEQ AGUARDA_CM	#Desvia se igual a 0 (botão não foi pressionado)
tmp(386) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(387) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(388) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do acumulador em MEM[15] (inibir centena de milhar)
tmp(389) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(390) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do acumulador no LDR9
tmp(391) := "00" & x"A" & '0' & x"00";	-- RET
tmp(392) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega 0 para o acumulador
tmp(393) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(394) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador na MEM[9] (flag inibir contagem)
tmp(395) := "00" & x"5" & '1' & x"FD";	-- STA 509, R0	#Limpa a leitura do botão KEY2
tmp(396) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	# Carrega MEM[0] (unidades) no acumulador
tmp(397) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[0] == 0
tmp(398) := "00" & x"7" & '1' & x"92";	-- JEQ VEMUM_D	# Se MEM[0] == 0, realiza o "empréstimo"
tmp(399) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[0]
tmp(400) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	# Armazena o novo valor de MEM[0]
tmp(401) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(402) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(403) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	# Define MEM[0] para 9
tmp(404) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	# Carrega MEM[1] (dezenas) no acumulador
tmp(405) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[1] == 0
tmp(406) := "00" & x"7" & '1' & x"9A";	-- JEQ VEMUM_C	# Se MEM[1] == 0, realiza o próximo "empréstimo"
tmp(407) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[1]
tmp(408) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	# Armazena o novo valor de MEM[1]
tmp(409) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(410) := "00" & x"4" & '0' & x"06";	-- LDI 6, R0	# Carrega 6 no acumulador
tmp(411) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	# Define MEM[1] para 6
tmp(412) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	# Carrega MEM[2] (centenas) no acumulador
tmp(413) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[2] == 0
tmp(414) := "00" & x"7" & '1' & x"A2";	-- JEQ VEMUM_M	# Se MEM[2] == 0, realiza o próximo "empréstimo"
tmp(415) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[2]
tmp(416) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	# Armazena o novo valor de MEM[2]
tmp(417) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(418) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(419) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	# Define MEM[2] para 9
tmp(420) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	# Carrega MEM[3] (milhares) no acumulador
tmp(421) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[3] == 0
tmp(422) := "00" & x"7" & '1' & x"AA";	-- JEQ VEMUM_DM	# Se MEM[3] == 0, realiza o próximo "empréstimo"
tmp(423) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[3]
tmp(424) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	# Armazena o novo valor de MEM[3]
tmp(425) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(426) := "00" & x"4" & '0' & x"06";	-- LDI 6, R0	# Carrega 6 no acumulador
tmp(427) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	# Define MEM[3] para 6
tmp(428) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	# Carrega MEM[4] (dezenas de milhares) no acumulador
tmp(429) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[4] == 0
tmp(430) := "00" & x"7" & '1' & x"B2";	-- JEQ VEMUM_CM	# Se MEM[4] == 0, realiza o próximo "empréstimo"
tmp(431) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[4]
tmp(432) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	# Armazena o novo valor de MEM[4]
tmp(433) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(434) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(435) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	# Define MEM[4] para 9
tmp(436) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	# Carrega MEM[5] (centenas de milhares) no acumulador
tmp(437) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[5] == 0
tmp(438) := "00" & x"7" & '1' & x"BA";	-- JEQ ZERA_HEX	# Zera se for menos que 0
tmp(439) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[5]
tmp(440) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	# Armazena o novo valor de MEM[5]
tmp(441) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(442) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(443) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador na MEM[0] (unidades)
tmp(444) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador na MEM[1] (dezenas)
tmp(445) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador na MEM[2] (centenas)
tmp(446) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador na MEM[6] (milhar)
tmp(447) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador na MEM[7] (dezena de milhar)
tmp(448) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do acumulador na MEM[8] (centena de milhar)
tmp(449) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador na MEM[9] (flag inibir contagem)
tmp(450) := "00" & x"A" & '0' & x"00";	-- RET


        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;