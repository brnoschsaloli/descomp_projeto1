library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Operacao_ULA_2bits, habLeituraMEM, habEscritaMEM 
      -- Inicializa os endereços:
tmp(0) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(1) := "00" & x"5" & '1' & x"20";	-- STA 288, R0	#Armazena o valor do acumulador em HEX0
tmp(2) := "00" & x"5" & '1' & x"21";	-- STA 289, R0	#Armazena o valor do acumulador em HEX1
tmp(3) := "00" & x"5" & '1' & x"22";	-- STA 290, R0	#Armazena o valor do acumulador em HEX2
tmp(4) := "00" & x"5" & '1' & x"23";	-- STA 291, R0	#Armazena o valor do acumulador em HEX3
tmp(5) := "00" & x"5" & '1' & x"24";	-- STA 292, R0	#Armazena o valor do acumulador em HEX4
tmp(6) := "00" & x"5" & '1' & x"25";	-- STA 293, R0	#Armazena o valor do acumulador em HEX5
tmp(7) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(8) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(9) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(10) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(11) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do acumulador no LDR9
tmp(12) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(13) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(14) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador em MEM[0] (unidades)
tmp(15) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador em MEM[1] (dezenas)
tmp(16) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador em MEM[2] (centenas)
tmp(17) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador em MEM[6] (milhares)
tmp(18) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador em MEM[7] (dezenas de milhares)
tmp(19) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do acumulador em MEM[8] (centenas de milhares)
tmp(20) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador em MEM[9] (flag inibir contagem)
tmp(21) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega o acumulador com o valor 9
tmp(22) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do acumulador em MEM[10] (inibir unidade)
tmp(23) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do acumulador em MEM[11] (inibir dezena)
tmp(24) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do acumulador em MEM[12] (inibir centena)
tmp(25) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do acumulador em MEM[13] (inibir milhar)
tmp(26) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do acumulador em MEM[14] (inibir dezena de milhar)
tmp(27) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do acumulador em MEM[15] (inibir centena de milhar)
tmp(28) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(29) := "00" & x"5" & '1' & x"FF";	-- STA 511, R0	#Limpa a leitura do botão zero
tmp(30) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(31) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(32) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(33) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(34) := "11" & x"4" & '0' & x"03";	-- LDI 3, R3	#COLUNA 3
tmp(35) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(36) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(37) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(38) := "11" & x"4" & '0' & x"12";	-- LDI 18, R3	#R
tmp(39) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(40) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(41) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#COLUNA 4
tmp(42) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(43) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(44) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(45) := "11" & x"4" & '0' & x"05";	-- LDI 5, R3	#E
tmp(46) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(47) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(48) := "11" & x"4" & '0' & x"05";	-- LDI 5, R3	#COLUNA 5
tmp(49) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(50) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(51) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(52) := "11" & x"4" & '0' & x"0C";	-- LDI 12, R3	#L
tmp(53) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(54) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(55) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#COLUNA 6
tmp(56) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(57) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(58) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(59) := "11" & x"4" & '0' & x"0F";	-- LDI 15, R3	#O
tmp(60) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(61) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(62) := "11" & x"4" & '0' & x"07";	-- LDI 7, R3	#COLUNA 7
tmp(63) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(64) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(65) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(66) := "11" & x"4" & '0' & x"07";	-- LDI 7, R3	#G
tmp(67) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(68) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(69) := "11" & x"4" & '0' & x"08";	-- LDI 8, R3	#COLUNA 8
tmp(70) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(71) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(72) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(73) := "11" & x"4" & '0' & x"09";	-- LDI 9, R3	#I
tmp(74) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(75) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(76) := "11" & x"4" & '0' & x"09";	-- LDI 9, R3	#COLUNA 9
tmp(77) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(78) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(79) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(80) := "11" & x"4" & '0' & x"0F";	-- LDI 15, R3	#O
tmp(81) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(82) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(83) := "11" & x"4" & '0' & x"0B";	-- LDI 11, R3	#COLUNA 11
tmp(84) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(85) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(86) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(87) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#B
tmp(88) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(89) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(90) := "11" & x"4" & '0' & x"0C";	-- LDI 12, R3	#COLUNA 12
tmp(91) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(92) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(93) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(94) := "11" & x"4" & '0' & x"01";	-- LDI 1, R3	#A
tmp(95) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(96) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(97) := "11" & x"4" & '0' & x"0D";	-- LDI 13, R3	#COLUNA 13
tmp(98) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(99) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(100) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(101) := "11" & x"4" & '0' & x"03";	-- LDI 3, R3	#C
tmp(102) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(103) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(104) := "11" & x"4" & '0' & x"0E";	-- LDI 14, R3	#COLUNA 14
tmp(105) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(106) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(107) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(108) := "11" & x"4" & '0' & x"01";	-- LDI 1, R3	#A
tmp(109) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(110) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(111) := "11" & x"4" & '0' & x"0F";	-- LDI 15, R3	#COLUNA 15
tmp(112) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(113) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(114) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(115) := "11" & x"4" & '0' & x"0E";	-- LDI 14, R3	#N
tmp(116) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(117) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(118) := "11" & x"4" & '0' & x"10";	-- LDI 16, R3	#COLUNA 16
tmp(119) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(120) := "11" & x"4" & '0' & x"02";	-- LDI 2, R3	#LINHA 2
tmp(121) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(122) := "11" & x"4" & '0' & x"01";	-- LDI 1, R3	#A
tmp(123) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(124) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(125) := "11" & x"4" & '0' & x"06";	-- LDI 6, R3	#COLUNA 6
tmp(126) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(127) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(128) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(129) := "11" & x"4" & '0' & x"30";	-- LDI 48, R3	#0
tmp(130) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(131) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(132) := "11" & x"4" & '0' & x"07";	-- LDI 7, R3	#COLUNA 7
tmp(133) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(134) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(135) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(136) := "11" & x"4" & '0' & x"30";	-- LDI 48, R3	#0
tmp(137) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(138) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(139) := "11" & x"4" & '0' & x"08";	-- LDI 8, R3	#COLUNA 8
tmp(140) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(141) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(142) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(143) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(144) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(145) := "11" & x"4" & '0' & x"09";	-- LDI 9, R3	#COLUNA 9
tmp(146) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(147) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(148) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(149) := "11" & x"4" & '0' & x"30";	-- LDI 48, R3	#0
tmp(150) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(151) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(152) := "11" & x"4" & '0' & x"0A";	-- LDI 10, R3	#COLUNA 10
tmp(153) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(154) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(155) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(156) := "11" & x"4" & '0' & x"30";	-- LDI 48, R3	#0
tmp(157) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(158) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(159) := "11" & x"4" & '0' & x"0B";	-- LDI 11, R3	#COLUNA 11
tmp(160) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(161) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(162) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(163) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(164) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(165) := "11" & x"4" & '0' & x"0C";	-- LDI 12, R3	#COLUNA 12
tmp(166) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(167) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(168) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(169) := "11" & x"4" & '0' & x"30";	-- LDI 48, R3	#0
tmp(170) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(171) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(172) := "11" & x"4" & '0' & x"0D";	-- LDI 13, R3	#COLUNA 13
tmp(173) := "11" & x"5" & '1' & x"80";	-- STA 384, R3	#ARMAZENA NO REGISTRADOR DAS COLUNAS
tmp(174) := "11" & x"4" & '0' & x"04";	-- LDI 4, R3	#LINHA 4
tmp(175) := "11" & x"5" & '1' & x"81";	-- STA 385, R3	#ARMAZENA NO REGISTRADOR DAS LINHAS
tmp(176) := "11" & x"4" & '0' & x"30";	-- LDI 48, R3	#0
tmp(177) := "11" & x"5" & '1' & x"82";	-- STA 386, R3	#ARMAZENA NO REGISTRADOR DA DATA
tmp(178) := "11" & x"5" & '1' & x"83";	-- STA 387, R3	#MANDA PRA VGA
tmp(179) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(180) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(181) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(182) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(183) := "00" & x"1" & '1' & x"60";	-- LDA 352, R0	#Carrega o acumulador com a leitura do botão KEY0
tmp(184) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(185) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(186) := "00" & x"7" & '0' & x"BD";	-- JEQ NAO_CLICOU0	#Desvia se igual a 0 (botão não foi pressionado)
tmp(187) := "00" & x"9" & '0' & x"D5";	-- JSR INCREMENTO	#O botão foi pressionado, chama a sub-rotina de incremento
tmp(188) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de incremento
tmp(189) := "00" & x"9" & '1' & x"0E";	-- JSR SALVA_DISP	#Escreve o valor das váriaveis de contagem nos displays
tmp(190) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de salvar nos displays
tmp(191) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(192) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(193) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(194) := "00" & x"7" & '0' & x"C5";	-- JEQ NAO_CLICOU1	#Desvia se igual a 0 (botão não foi pressionado)
tmp(195) := "00" & x"9" & '1' & x"48";	-- JSR DEFINE_LIM	#O botão foi pressionado, chama a sub-rotina de incremento
tmp(196) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de definir limite
tmp(197) := "00" & x"9" & '1' & x"2C";	-- JSR VERIFICA_LIM
tmp(198) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de verificar limite
tmp(199) := "00" & x"1" & '1' & x"62";	-- LDA 354, R0	#Carrega o acumulador com a leitura do botão KEY2
tmp(200) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(201) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(202) := "00" & x"7" & '0' & x"CD";	-- JEQ NAO_CLICOU2	#Desvia se igual a 0 (botão não foi pressionado)
tmp(203) := "00" & x"9" & '1' & x"7D";	-- JSR DECREMENTO	#O botão foi pressionado, chama a sub-rotina de incremento
tmp(204) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de incremento
tmp(205) := "00" & x"1" & '1' & x"64";	-- LDA 356, R0	#Carrega o acumulador com a leitura do botão FPGA_RESET
tmp(206) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(207) := "00" & x"D" & '0' & x"01";	-- CEQi 1, R0	#Compara com constante 1
tmp(208) := "00" & x"7" & '0' & x"D2";	-- JEQ REINICIO	#Desvia se igual a 1 (botão não foi pressionado)
tmp(209) := "00" & x"9" & '1' & x"1B";	-- JSR RESET	#O botão foi pressionado, chama a sub-rotina de reset
tmp(210) := "00" & x"0" & '0' & x"00";	-- NOP	#Retorno da sub-rotina de reset
tmp(211) := "00" & x"6" & '0' & x"B6";	-- JMP INICIO	#Fecha o laço principal, faz uma nova leitura de KEY0
tmp(212) := "00" & x"0" & '0' & x"00";	-- NOP
tmp(213) := "00" & x"5" & '1' & x"FF";	-- STA 511, R0	#Limpa a leitura do botão
tmp(214) := "00" & x"1" & '0' & x"09";	-- LDA 9, R0	#Carrega o valor de MEM[9] (flag inibir contagem)
tmp(215) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara o valor com constante 0
tmp(216) := "00" & x"7" & '0' & x"DA";	-- JEQ INCREMENTAR
tmp(217) := "00" & x"A" & '0' & x"00";	-- RET
tmp(218) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	#Carrega o valor de MEM[0] (contador)
tmp(219) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(220) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(221) := "00" & x"7" & '0' & x"E0";	-- JEQ VAIUM_D	#Realiza o carry out caso valor igual a 10
tmp(222) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Salva o incremento em MEM[0] (contador)
tmp(223) := "00" & x"A" & '0' & x"00";	-- RET	#Retorna da sub-rotina
tmp(224) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(225) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador em MEM[0] (unidades)
tmp(226) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	#Carrega valor de MEM[1] no acumulador (dezenas)
tmp(227) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(228) := "00" & x"D" & '0' & x"06";	-- CEQi 6, R0	#Compara o valor com constante 10
tmp(229) := "00" & x"7" & '0' & x"E8";	-- JEQ VAIUM_C	#Realiza o carry out caso valor igual a 10
tmp(230) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Salva o incremento em MEM[1] (dezenas)
tmp(231) := "00" & x"A" & '0' & x"00";	-- RET
tmp(232) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(233) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador em MEM[1] (dezenas)
tmp(234) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	#Carrega valor de MEM[2] no acumulador (centenas)
tmp(235) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(236) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(237) := "00" & x"7" & '0' & x"F0";	-- JEQ VAIUM_M	#Realiza o carry out caso valor igual a 10
tmp(238) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Salva o incremento em MEM[2] (centenas)
tmp(239) := "00" & x"A" & '0' & x"00";	-- RET
tmp(240) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(241) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador em MEM[2] (centenas)
tmp(242) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	#Carrega valor de MEM[6] no acumulador (milhares)
tmp(243) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(244) := "00" & x"D" & '0' & x"06";	-- CEQi 6, R0	#Compara o valor com constante 10
tmp(245) := "00" & x"7" & '0' & x"F8";	-- JEQ VAIUM_DM	#Realiza o carry out caso valor igual a 10
tmp(246) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Salva o incremento em MEM[6] (milhares)
tmp(247) := "00" & x"A" & '0' & x"00";	-- RET
tmp(248) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(249) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador em MEM[6] (milhares)
tmp(250) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	#Carrega valor de MEM[7] no acumulador (dezenas de milhares)
tmp(251) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(252) := "01" & x"1" & '0' & x"08";	-- LDA 8, R1	#Carrega valor de MEM[8] no acumulador (centenas de milhares)
tmp(253) := "01" & x"D" & '0' & x"02";	-- CEQi 2, R1	#Compara o valor com constante 2
tmp(254) := "00" & x"7" & '1' & x"02";	-- JEQ COMPARA4	#Pula para o fim da rotina
tmp(255) := "00" & x"D" & '0' & x"0A";	-- CEQi 10, R0	#Compara o valor com constante 10
tmp(256) := "00" & x"7" & '1' & x"06";	-- JEQ VAIUM_CM	#Realiza o carry out caso valor igual a 10
tmp(257) := "00" & x"6" & '1' & x"04";	-- JMP END_DM
tmp(258) := "00" & x"D" & '0' & x"04";	-- CEQi 4, R0	#Compara o valor com constante 4
tmp(259) := "00" & x"7" & '1' & x"06";	-- JEQ VAIUM_CM	#Realiza o carry out caso valor igual a 4
tmp(260) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Salva o incremento em MEM[7] (dezenas de milhares)
tmp(261) := "00" & x"A" & '0' & x"00";	-- RET
tmp(262) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega valor 0 no acumulador (constante 0)
tmp(263) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador em MEM[7] (dezenas milhares)
tmp(264) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega valor de MEM[8] no acumulador (centenas de milhares)
tmp(265) := "00" & x"E" & '0' & x"01";	-- ADDi 1, R0	#ADDi com a constante 1
tmp(266) := "00" & x"D" & '0' & x"03";	-- CEQi 3, R0	#Compara o valor com constante 3
tmp(267) := "00" & x"7" & '1' & x"AF";	-- JEQ ZERA_HEX	#Zera se chegar ao final
tmp(268) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Salva o incremento em MEM[8] (centena de milhares)
tmp(269) := "00" & x"A" & '0' & x"00";	-- RET
tmp(270) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	#Carrega o valor de MEM[0] (unidades)
tmp(271) := "00" & x"5" & '1' & x"20";	-- STA 288, R0	#Armazena valor do acumulador de unidades no HEX0
tmp(272) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	#Carrega o valor de MEM[1] (dezenas)
tmp(273) := "00" & x"5" & '1' & x"21";	-- STA 289, R0	#Armazena valor do acumulador de dezenas no HEX1
tmp(274) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	#Carrega o valor de MEM[2] (centenas)
tmp(275) := "00" & x"5" & '1' & x"22";	-- STA 290, R0	#Armazena valor do acumulador de centenas no HEX2
tmp(276) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	#Carrega o valor de MEM[6] (milhares)
tmp(277) := "00" & x"5" & '1' & x"23";	-- STA 291, R0	#Armazena valor do acumulador de unidades no HEX3
tmp(278) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	#Carrega o valor de MEM[7] (dezenas de milhares)
tmp(279) := "00" & x"5" & '1' & x"24";	-- STA 292, R0	#Armazena valor do acumulador de dezenas no HEX4
tmp(280) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega o valor de MEM[8] (centenas de milhares)
tmp(281) := "00" & x"5" & '1' & x"25";	-- STA 293, R0	#Armazena valor do acumulador de centenas no HEX5
tmp(282) := "00" & x"A" & '0' & x"00";	-- RET
tmp(283) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(284) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador na MEM[0] (unidades)
tmp(285) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador na MEM[1] (dezenas)
tmp(286) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador na MEM[2] (centenas)
tmp(287) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador na MEM[6] (milhar)
tmp(288) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador na MEM[7] (dezena de milhar)
tmp(289) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do acumulador na MEM[8] (centena de milhar)
tmp(290) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador na MEM[9] (flag inibir contagem)
tmp(291) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(292) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	#Carrega o acumulador com o valor 9
tmp(293) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do acumulador em MEM[10] (inibir unidade)
tmp(294) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do acumulador em MEM[11] (inibir dezena)
tmp(295) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do acumulador em MEM[12] (inibir centena)
tmp(296) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do acumulador em MEM[13] (inibir milhar)
tmp(297) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do acumulador em MEM[14] (inibir dezena de milhar)
tmp(298) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do acumulador em MEM[15] (inibir centena de milhar)
tmp(299) := "00" & x"A" & '0' & x"00";	-- RET
tmp(300) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	#Carrega o valor de MEM[0] (unidades)
tmp(301) := "00" & x"8" & '0' & x"0A";	-- CEQ 10, R0	#Compara o valor de MEM[10] (inibir unidade)
tmp(302) := "00" & x"7" & '1' & x"30";	-- JEQ NEXT_LIM1
tmp(303) := "00" & x"A" & '0' & x"00";	-- RET
tmp(304) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	#Carrega o valor de MEM[1] (dezenas)
tmp(305) := "00" & x"8" & '0' & x"0B";	-- CEQ 11, R0	#Compara o valor de MEM[11] (inibir dezenas)
tmp(306) := "00" & x"7" & '1' & x"34";	-- JEQ NEXT_LIM2
tmp(307) := "00" & x"A" & '0' & x"00";	-- RET
tmp(308) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	#Carrega o valor de MEM[2] (centenas)
tmp(309) := "00" & x"8" & '0' & x"0C";	-- CEQ 12, R0	#Compara o valor de MEM[12] (inibir centenas)
tmp(310) := "00" & x"7" & '1' & x"38";	-- JEQ NEXT_LIM3
tmp(311) := "00" & x"A" & '0' & x"00";	-- RET
tmp(312) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	#Carrega o valor de MEM[6] (milhar)
tmp(313) := "00" & x"8" & '0' & x"0D";	-- CEQ 13, R0	#Compara o valor de MEM[13] (inibir milhar)
tmp(314) := "00" & x"7" & '1' & x"3C";	-- JEQ NEXT_LIM4
tmp(315) := "00" & x"A" & '0' & x"00";	-- RET
tmp(316) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	#Carrega o valor de MEM[7] (dezena de milhar)
tmp(317) := "00" & x"8" & '0' & x"0E";	-- CEQ 14, R0	#Compara o valor de MEM[10] (inibir dezena de milhar)
tmp(318) := "00" & x"7" & '1' & x"40";	-- JEQ NEXT_LIM5
tmp(319) := "00" & x"A" & '0' & x"00";	-- RET
tmp(320) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	#Carrega o valor de MEM[8] (centena de milhar)
tmp(321) := "00" & x"8" & '0' & x"0F";	-- CEQ 15, R0	#Compara o valor de MEM[10] (inibir centena de milhar)
tmp(322) := "00" & x"7" & '1' & x"44";	-- JEQ TODOS_IGUAL
tmp(323) := "00" & x"A" & '0' & x"00";	-- RET
tmp(324) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o acumulador com o valor 1
tmp(325) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador em MEM[9] (flag inibir contagem)
tmp(326) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(327) := "00" & x"A" & '0' & x"00";	-- RET
tmp(328) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(329) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(330) := "00" & x"5" & '0' & x"0A";	-- STA 10, R0	#Armazena o valor do acumulador em MEM[10] (inibir unidade)
tmp(331) := "00" & x"4" & '0' & x"04";	-- LDI 4, R0	#Carrega o acumulador com o valor 4
tmp(332) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(333) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(334) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(335) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(336) := "00" & x"7" & '1' & x"4D";	-- JEQ AGUARDA_D	#Desvia se igual a 0 (botão não foi pressionado)
tmp(337) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(338) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(339) := "00" & x"5" & '0' & x"0B";	-- STA 11, R0	#Armazena o valor do acumulador em MEM[11] (inibir dezena)
tmp(340) := "00" & x"4" & '0' & x"10";	-- LDI 16, R0	#Carrega o acumulador com o valor 16
tmp(341) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(342) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(343) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(344) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(345) := "00" & x"7" & '1' & x"56";	-- JEQ AGUARDA_C	#Desvia se igual a 0 (botão não foi pressionado)
tmp(346) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(347) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(348) := "00" & x"5" & '0' & x"0C";	-- STA 12, R0	#Armazena o valor do acumulador em MEM[12] (inibir centena)
tmp(349) := "00" & x"4" & '0' & x"20";	-- LDI 32, R0	#Carrega o acumulador com o valor 32
tmp(350) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(351) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(352) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(353) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(354) := "00" & x"7" & '1' & x"5F";	-- JEQ AGUARDA_M	#Desvia se igual a 0 (botão não foi pressionado)
tmp(355) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(356) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(357) := "00" & x"5" & '0' & x"0D";	-- STA 13, R0	#Armazena o valor do acumulador em MEM[13] (inibir milhar)
tmp(358) := "00" & x"4" & '0' & x"80";	-- LDI 128, R0	#Carrega o acumulador com o valor 128
tmp(359) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(360) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(361) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(362) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(363) := "00" & x"7" & '1' & x"68";	-- JEQ AGUARDA_DM	#Desvia se igual a 0 (botão não foi pressionado)
tmp(364) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(365) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(366) := "00" & x"5" & '0' & x"0E";	-- STA 14, R0	#Armazena o valor do acumulador em MEM[13] (inibir dezena de milhar)
tmp(367) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(368) := "00" & x"5" & '1' & x"00";	-- STA 256, R0	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(369) := "00" & x"4" & '0' & x"01";	-- LDI 1, R0	#Carrega o acumulador com o valor 1
tmp(370) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do acumulador no LDR9
tmp(371) := "00" & x"1" & '1' & x"61";	-- LDA 353, R0	#Carrega o acumulador com a leitura do botão KEY1
tmp(372) := "00" & x"C" & '0' & x"01";	-- ANDi 1, R0	#Utiliza a máscara b0000_0001 para limpar todos os bits menos o bit 0
tmp(373) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	#Compara com constante 0
tmp(374) := "00" & x"7" & '1' & x"73";	-- JEQ AGUARDA_CM	#Desvia se igual a 0 (botão não foi pressionado)
tmp(375) := "00" & x"5" & '1' & x"FE";	-- STA 510, R0	#Limpa a leitura do botão um
tmp(376) := "00" & x"1" & '1' & x"40";	-- LDA 320, R0	#Carrega o acumulador com a leitura do SW7TO0
tmp(377) := "00" & x"5" & '0' & x"0F";	-- STA 15, R0	#Armazena o valor do acumulador em MEM[15] (inibir centena de milhar)
tmp(378) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(379) := "00" & x"5" & '1' & x"02";	-- STA 258, R0	#Armazena o valor do bit0 do acumulador no LDR9
tmp(380) := "00" & x"A" & '0' & x"00";	-- RET
tmp(381) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega 0 para o acumulador
tmp(382) := "00" & x"5" & '1' & x"01";	-- STA 257, R0	#Armazena o valor do bit0 do acumulador no LDR8
tmp(383) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador na MEM[9] (flag inibir contagem)
tmp(384) := "00" & x"5" & '1' & x"FD";	-- STA 509, R0	#Limpa a leitura do botão KEY2
tmp(385) := "00" & x"1" & '0' & x"00";	-- LDA 0, R0	# Carrega MEM[0] (unidades) no acumulador
tmp(386) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[0] == 0
tmp(387) := "00" & x"7" & '1' & x"87";	-- JEQ VEMUM_D	# Se MEM[0] == 0, realiza o "empréstimo"
tmp(388) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[0]
tmp(389) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	# Armazena o novo valor de MEM[0]
tmp(390) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(391) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(392) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	# Define MEM[0] para 9
tmp(393) := "00" & x"1" & '0' & x"01";	-- LDA 1, R0	# Carrega MEM[1] (dezenas) no acumulador
tmp(394) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[1] == 0
tmp(395) := "00" & x"7" & '1' & x"8F";	-- JEQ VEMUM_C	# Se MEM[1] == 0, realiza o próximo "empréstimo"
tmp(396) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[1]
tmp(397) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	# Armazena o novo valor de MEM[1]
tmp(398) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(399) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(400) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	# Define MEM[1] para 9
tmp(401) := "00" & x"1" & '0' & x"02";	-- LDA 2, R0	# Carrega MEM[2] (centenas) no acumulador
tmp(402) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[2] == 0
tmp(403) := "00" & x"7" & '1' & x"97";	-- JEQ VEMUM_M	# Se MEM[2] == 0, realiza o próximo "empréstimo"
tmp(404) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[2]
tmp(405) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	# Armazena o novo valor de MEM[2]
tmp(406) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(407) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(408) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	# Define MEM[2] para 9
tmp(409) := "00" & x"1" & '0' & x"06";	-- LDA 6, R0	# Carrega MEM[3] (milhares) no acumulador
tmp(410) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[3] == 0
tmp(411) := "00" & x"7" & '1' & x"9F";	-- JEQ VEMUM_DM	# Se MEM[3] == 0, realiza o próximo "empréstimo"
tmp(412) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[3]
tmp(413) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	# Armazena o novo valor de MEM[3]
tmp(414) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(415) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(416) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	# Define MEM[3] para 9
tmp(417) := "00" & x"1" & '0' & x"07";	-- LDA 7, R0	# Carrega MEM[4] (dezenas de milhares) no acumulador
tmp(418) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[4] == 0
tmp(419) := "00" & x"7" & '1' & x"A7";	-- JEQ VEMUM_CM	# Se MEM[4] == 0, realiza o próximo "empréstimo"
tmp(420) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[4]
tmp(421) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	# Armazena o novo valor de MEM[4]
tmp(422) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(423) := "00" & x"4" & '0' & x"09";	-- LDI 9, R0	# Carrega 9 no acumulador
tmp(424) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	# Define MEM[4] para 9
tmp(425) := "00" & x"1" & '0' & x"08";	-- LDA 8, R0	# Carrega MEM[5] (centenas de milhares) no acumulador
tmp(426) := "00" & x"D" & '0' & x"00";	-- CEQi 0, R0	# Verifica se MEM[5] == 0
tmp(427) := "00" & x"7" & '1' & x"AF";	-- JEQ ZERA_HEX	# Zera se for menos que 0
tmp(428) := "00" & x"F" & '0' & x"01";	-- SUBi 1, R0	# Subtrai 1 de MEM[5]
tmp(429) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	# Armazena o novo valor de MEM[5]
tmp(430) := "00" & x"A" & '0' & x"00";	-- RET	# Retorna da sub-rotina
tmp(431) := "00" & x"4" & '0' & x"00";	-- LDI 0, R0	#Carrega o acumulador com o valor 0
tmp(432) := "00" & x"5" & '0' & x"00";	-- STA 0, R0	#Armazena o valor do acumulador na MEM[0] (unidades)
tmp(433) := "00" & x"5" & '0' & x"01";	-- STA 1, R0	#Armazena o valor do acumulador na MEM[1] (dezenas)
tmp(434) := "00" & x"5" & '0' & x"02";	-- STA 2, R0	#Armazena o valor do acumulador na MEM[2] (centenas)
tmp(435) := "00" & x"5" & '0' & x"06";	-- STA 6, R0	#Armazena o valor do acumulador na MEM[6] (milhar)
tmp(436) := "00" & x"5" & '0' & x"07";	-- STA 7, R0	#Armazena o valor do acumulador na MEM[7] (dezena de milhar)
tmp(437) := "00" & x"5" & '0' & x"08";	-- STA 8, R0	#Armazena o valor do acumulador na MEM[8] (centena de milhar)
tmp(438) := "00" & x"5" & '0' & x"09";	-- STA 9, R0	#Armazena o valor do acumulador na MEM[9] (flag inibir contagem)
tmp(439) := "00" & x"A" & '0' & x"00";	-- RET


        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;